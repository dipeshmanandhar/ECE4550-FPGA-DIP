��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����A�
&CʁRR���o>���q+�AR��k�b� B�����C(D�x)�d�!gN&{����+&f���^��T�JЬJ	yh�ldڪ��:RV۽�أv��椏"�c!����2���I�U<�? 5p��ݩ�L=L�E
�N�`^Ӿ��$Zϩ_�-�,S4��,�Wl�Sņ�4tr}(.`<3�e���ݍ�A���M��2�n"��\�t�H�&� ��z�~rfяܞ}�7� ��fUiҝ������l3��oTq%���B"u�� Ej��F��Y�ԸJJ4
���[���.�����9��S��M[����� ��J)���wB+�j�IBfiҁ7GLR�QxU�'��N-��%��Ѝl�q�2���6�}L�݂h�l���k3/ro�f�[����]?pƒF�R_��]�a��Y�5�)��%}1��0bɞ&���m_�����F$�w�����o��%��2LOB��ܰ���i��)$e��t�Ⱦ�`�84�Bp�P����q�@�z7��Mɻ���1��M����@�����l�!/�Q�\����Y�x���D�/�����G�}��4af���.BP�ʽ�!�r	9����I���'=���j�Uk ���BF���R��Y�����zZr���r���O�Ui��|o����I��U,/Dbf+� ���&1۫��Y;���6��iQ���!C�覊��Mж	H��<j*���LZ�(�#؁ ���c�[�0t���6h�Q�H�~�T؀Ǎ�J� ��_{���H�]Ð�$�R6�[����D �m2�TZJ�B1�>	��<�q����j�$ۏF�J���������Q`�hiJ��S*NqKx�e6�O�?"|.š�k���O�8lWB���'a8�YY�ʆZKаϡG�c�8p�PGE�eaE���=?)J�.!,��=Ŀ�q�LJ�����Q9�BTm�]��suZWA���On��C�v�!�~����&��ر�OL]G�Y˽1���
��tY�(��h8���4>��F�F��_�\��~��!&Z�]�	�F�fz?��{o���z�BJ �ߧ�� 9����f\���?K	z��Qr�;��w1*��`��JARAY6���ܝR���.o�1Z��d[�*�&�6�c*�8�B%��E�x�I��ưf�r�+��1z��cS�D>�Dc��H�ŋ�/c��@Ҷ>���^r{�Y��b�!�F�B�-e"����7��aХˬٞ�� 7�� 6 �Y�D{��~�>{E���~f �]�"��{dB2�o�Jl��O ~B���&�t��g�h����{5�K�r4�_y%HU?��!�n�� fa��֞�� �����>L)4�enZ޾:�K�������㳀�pYbG����ʆ	&�-�1�$����:ؕb��l#"���^Z�`Z������}B(�&�m/m�|���K<�
�8�> �k�g��Վy�r<�ApC���T�J�"�:��x���|F�q+Ɋ�DY��4'�s�E1\�y�����Q��w�@�SJW����\���*�[%�4��8m6&�Fy�ޱu�胈������ᡧ�z���Tl�ZY�!j�NT�`��[��r�G踓����'�{�"�0i�i�t��4zSԤ�5���)]ؿ��֋�킐$���9�,�9́m1v�*��l>���h�^���Ú���~՚��|p�E�ą^C�Ԫc�y�噭��!��%����f��A�����ɰA!��[�a�LFF�_ɔ����*1��!��caOэbz�o9��(O�}W�t�N�@Z�I<���%:���T�y�]5Z�W ܭ�SGwU��4j\�nze����}R��f�%��x������+epKuih&�H�����P�VȎ٘1��s�u�,_������q�o'.��Gj(��. �y�^~9�w� ��ѱѩ='L�:�c0��Z�x�WD����z>���s��`�&*1�5]&p+,b�.zr�����֟!n�}X��Z,䷇�Z��S ��_ynT�Ck���'�R��v���a��i��l��?j&d��G��<� �_L)F���C^۰P��-����-�Fs��ِZm\���Gֿ�7��),o{�3X7������@��O-��G�˲����	�1Y$M��*)\XL�aB�����dY.����=�wF�!�����8$^�Aw,;�5����N{C�>o0���-r��e���34�˟{(����jD��ܵ�e���k��'�l��l2�5���|X7W�ѯT�PP������ʛn$ec7v���r ��>e=, Ĩ�䨧�+�#<ܓ�L�O�'!o�-O3�\�>j������g�S̩olns�_�'���g�����m���������CQ��o���r��,���b��i����;Tm�fA��"J���Q�N�Б����@�~��h�Β&�QB/���?C�p�jۀ&�]*�ד-��8�^�U�R�>̣��"nC���'�����vɥ�_��}�cL��5kTȚ4Ջ��J�a�ZǕ7���_R��Au�H/]�����Tz؟�&�����#�V����+�<�h�����SJ��0��^�J;�TRs�	����#�Œn�zXFNi�+WϑG�HG���+��a S������e �L��[����3i��?s�BU�F̙(�Oq�4�~{#� �c�ɠG���#��8�MP�Y���C��*"�R����KQ8�̗����|7��z3�+�)�Q'�K�['��.i�=��(�m�Z9���)0d~���	��[�������<%07�_��!��Q��d9�g�BU#R��ez��T8�T���w8@�lۀD�0wʞ��,P�;Ś��R"@c�`Ci�6��ue�� ��N�~q<��GC.0T��۹�Ʃ�T���R��ca�v�p8�l����"�᝺�J�kJ��i[��f�	l�bi=���r�}2r���kzI�>��ky6w̸����c��"���MC�`�ݝQ�����JS�������3��ߑ8Ds"�����/Y�}2����rO������{�kذ��p۽ߣ\��>��sdh�(gx��&w0�Ԟ� ����b**���B9���_������:�@��AMQ����9�DZE��,1�$��N�V ��7�tZx�ә�9��qZ��ЄF�"��[�߬���fQ�BFּo��v9�1ϋ���X�k�1p(�Z�E�MNj�(li����c���i������Vx��o�g*	u0՜�dG�q����G�aq�L�_���V\���!�)����;,�-���D�9��>�/.�--�OrMN�¸�أ�i�o��Ɵ�17���빾t���$��e&�'!����xm���*j�.��5��֋Ƚ�}��ae��H{Yz�0��I�M&X�"N�ݸ�ŶŞ�ב�5�?;�m�QQR��̄�)ЧCc�0�"CM����]��(=pz� A�.��<�q�k�຀��r����j����Z����'��;�$P�5V哅9RF�)m`�7�V�݉닩���ص
F�{�ͫ$7���T q}Ա�?���'��E&�%;�˝����d��A��Ӫ7��۫�Z��]W�~ʵy�8]QH�'uF5�IV<�K�t��R�({>����0Q��!<j!��4YzFh��´z��^��}oZp���&�X]hF�r7]��8{b���uK���QmB�@�O��jB�K�����/�\�nAs�	V�_�ٔ ⡉�:&�T�ߠ��!��? lP)�L����3��ZR���f�;��� 4 	��)IM�4㢯�Ps��0��'�`Ɯ�`EH�.�C��K��䏁���`�8R�9{��^����u�?��p�+Of������3li>�Lgg�����6�������z�'U"jn��<�6� 4�	8X�;�Z�:�àۤٗ��S"�7�'�p)$���!�X��wo[��F����X�+e�7�:�l�=��Y-����R;��?���-+����ĵ}�27;;�����j���4���;��2��x"��ܵ*%ŚX�� <�/;�Ӣ��I��Q��/׺+�A�����}�(�(b���Ԓu��iZ����e.��%���y>�C���R1�a6VX�������ɑ�F95�>��{��([���\\\� ��mW@�a�Zbܲ
�����/�.ܞ)�p+����h���M2��9�3PqU�`cq@Rp|�-*D}�a¢<����3ԋ���~�U���ls
�r��g��կ�ĩQ2xkt�������*���]�q�`�:A��o��Y��@����W��NZ�<{��
:X�ݲ����C�Ozs�}lLU���+��Oޯ
y�3�y֭�#D�}~���"�ďX��1nG� ��V2�eSxξ;�N���)���ܿ���(;��8��#��	*���f	ےD�rnI2x)9{�pݟ?�D5�63�#���:�
�RNK�So�&�j@�O�/V>��ȸN
OY��b�4F%K�蜅��d��j?樿P�Q.��u�Ͳ�d|�N`}��Z��A�In�[�lM^%P;NM�����f��!l���\�Z�XWm[�S����C.w�M�@'.�$�Z��W[>��ɚB�,(��R*I-�ܟ��)�\m������[�Sc8Ab�$�H�wdMJCE�ć������ן�k<�;/���+�H5O�I�E��������#
|_��D�eT7����a�ݛ^o�QwtΝ*O���t�Hs[�޴���n���Nc�'ձ�r�D�n�������g���Z *���H���/]��)�;��]�ӏ���ƙ�@V�Ӌ��|�s\/�&���)����i~��f��LHky�#^fl]5�#��i)@5W��Câu��
�#.��"��.n��-���s�Y�z!�rGIK���4Ѽ�Ns����c���E |[�0!�������tT���{������M�1ݬ��6�]6�!�A�<x_����F��u1Wk>�;��c�D埤P��C`���h��F��_h�2�r{��ŦK�=�~�	8�~�joڦ�&�K�q�ǿ��n�N�.=�Wl���ϖ��~Z�˕D��M~~�����֗����_�u���	��Tn��5k����<H�2p�V��l0O�3�����#���x-�����E'����%'��67��� "���#���ou��A�Yꯜ6���V���>F3洅�u��-z�R�2.`X�&����� >�+�'�F���M�#P��K�0j��qQ앢��6�0U,��}d���&�y�d�Q@�N�3��,���zU�c�M�bz�9��@����ܠ��]�D��.��p|u��i$�{wf�	��q�M�`��G�����˕��oVJ��jYvU��7ar�� ��Cv��}�i��M���/���r�2�@<�iH��C�5�/�抂�)����D�ח��7o��D�����򭨬Z/��e�U�|�>�@_�$���%8�y���`��u�B� �6t�+�PLrJi%)Ĩ�J��EpW�$�����2�5�	�����=#�L"��ڵY	��������:�Kїٵ�YKNj�j<IK�1T���^�8��to����w]��P]���Xϙp)��T<C�	����k��hC�{���Ba"��E��.�(��/L��ek�ikI�k�m?#'/�N�Qk�ͽ&Z�8�
����v���ę1d����#�J����n>\4v/�V�nGLsӔ��
�gm�0dK��:�U�o�\[rIןB��,��9��5�g�{��,����8�~1ӆK��~�i(��,;2�/2޺�~����M���&79�ľPB�j���Dok�K���7��C�CZfB��p�"G=��v�.;�,|�㎨�kV�>F�i�.3���f��D��ï���'[̝jH�=��+��ou�HԄļ��u�ߍN"=TS{����'�8)H��=A��](��
����l��/b+�<`-���b�|!�$�:&��4(�֐�S�9��p���5jFuv'�I�K� ����\DD�H������d��z?���=h���]f���~/x��lU�ZS�Ϝ�Q<z�ۧ�,`Ip�I'$T�s�K\o�����º�L�ן��}��ܘT�o>�7�[��8� ��a����l�3��7�ր#O�l��joi� e�����c�N�SLz�z�3��-9R�\���^�$��(֡�7jKZeko��q��������dD�ܬ�P	���զ�)=�ɞ6�
|H�Ku��)�	�
g`�<�+]���@I��y�̲~�w?�R߈���<l�>y���4s�-��p� Xkmӈ�9V�s���	�❱��e\���ɣx�j9#�.�gl�:/��6ռ��h(&BH�p%�;�����nՎ�zTk�w�f�#��hEe@d��lA���|�ݛJ]��%�SrC�Q��uK��ɟ���.{,�FieE%� ��w
�)3�[7e��	:�m}�IԶ�u���k��6��Ｏ�kJ�4O����~��齓8m?,I��Ğ���\������'�"�\N`Ov��ՋX�!j�;�O=n�
���iӟ�*yi�ʞ���v;���*I�ʳ�)�A�E����9c�t6�(V�--���OG�OZ-=۲1����)�J���'�/��wda�����)���oC��!��j>��k�YL�z�oI݉g����½%�@Q�j��\O��|<^ x)������t�X�8�,-�<2z��\#T�Q�u�P��ƻ�h��#etr�@��G1<d��8>�1��ah�/mt?v9?���O�&��"�cR�A�7ݧ�W�b-BJ�I��<?����W����Y�jn����-�+`�\ 5��|�g!$f���#~L&�t�c�q�j<����&eN��o��zG����B.+b	6_>�0�o�2H���h
�ä��
�K��J� �� �HFb(� ���aY�6��/��z~G)ԉ�2|��2�o�drl�e~E姽��]����ܡ�[�ohe��<���8~�Ut=XA�V_�T�<bi��������B�����)�J_����p�2_iDY�"�Ӷq��_R�8�@�Dz�v��
�~�Ȃx�aY�\ÐqG������C�C1���J1;�(L�3�E(] w�Z��a�t+y�<q���4�Z*�M��HU�޶�֦>�5:�y�w
h7��O��CH�b�]C:�P�ҝ`'mة$(ӪL��?ś��Gq�Ox����Z�u�ޝ�3ؖ����Q�_�=Xw[0��|�/��X�@<e5ԣg�p��N#�T4A�?agn' 3�-�0�GR&r�g���XS�Ɨ�i�m��SЧ����8]OґeFdʖr�	������D��xP�t3�/k����҂�f�=����o�I�DOY���тjoS4�Ɛ�%]�^5@�ux�nkt���R����'m�pQD�Կ\'0�<��o}/�m!bO�쿗�f͡r ��*O�Zv��Ӥ*ʰZ�n�:�c:1��,�$�*��p�Z���Kf�-_J7���GKe��Ps�<�cl+�5OY���:�Y�{=�qH�}�7��.f��rm�_w?�*���נh����d.���
kLN1�d|E��f���\`����n5�`G@��L�V�����k&@�pİ�=���J�=�l;	��|��/��2����I>K���θ�Ct��iE��%�vI&�q��]���9C��6sG�����̍>�1@Ch�>�Oݞ�̴�q<���-�P{�|����TigCl�/xoc&8���=�������& ��a�ى�y�	����պ%0rr��M�Y���0���emGxE�!����7E�tc=-�̝V�U_j?��!�[ ��	cx���Ȟ-bP� ��u���od9�F�����p7��KK�u�o���A��:Q��+C�e�Ϩ����ܣ��6q�Kxtl�6�8iޟ�U��I1��+6��T����L@ ��4�Ȩ~��ը��p�y�?��r��Z��=@J�����ϳ�Q�D� ;`��.Yv@Zx��B����;��SuE
:#v-4d��OO�Fy��5͖�Dv����|\�#��{L ��N���mB��&_R
6��_�ur�����Z�(����BW�i�!��/ET��De��wx&EIisP����7��`�>�k��I���z'=�Gly��3.�6M����P�%tm �Ju��¹B,�q���$�q]��^�i�� �$���)��VD:���*��gCh_ݢ�<�eԋ ��`}����@S�<�&�q6.�.�|�r��Ζo��wh��%T�[~~)o�eV�%�'E�c��"c�*(������N�:���ڰ�=c�x�OA�����FC�nT��DA�)��<�V:�@j��x��X:QBb��$�^s�����ɢuWN|�|�[L�y�.\PT��t����\�#��a�7 ���MBo�k�d�Pυy�ze$�<h&���vZ���Mq��2Բ|���O����9��8�k���
����X*"}���������Ug�ezb<��.Wȉ�:JfT��w(0vE�3�Ş����8
<	����aǈ��Ie��xE)�)Terw���Ⱥ!*m0���F��
Զ,���:����G8��	}�W����I��OA-�4�A�^�>z�� ��M������	�0�]D��Y�9k@e�w�ȳ��GTe�t�,#*pN�:�-�hun��<�	��բ)��*(���̻zV�Ѽ���%nЖд�5R�5)��x��j���%;���#4�*���8��[d�j=��ϙ�)���#u��|ſ��M%��b��FH�+��\X.�	�J1����YD�'����n3?��I�����"}A��u	5P����bV��b�i�c�:6/h�{��D��g���]��?��Ϛ�"ܽ�v2�6+j�G��,�NTR�L�$)��`8��a�d����9�����LcC1���S�GE^n ����u��x� ����^n�,N��eL_���Qņ�J�X?T�%t!���G Z�TS3���W ?��^H�]�������_Y37a�[:�m���"��OF{S��Y��J�mX�-j��e*8z�6b���f�/��?�jz��:�O����&t��o�"�E0�1�)�;v�����'CW�[�?|nW��U������߉�1T%7�=Q��_;��)�kz#�b���K��N��'Q���r���H�����q�>)	�������0
_fq��|{�l���'������Yv�����ĵ��ɞ�=�-o4�&�l���&�9�]4�����R\��9�L�O�ڊm�~3PQ�^�QjЪ`����e�S�$�n� ^��=�"r��2�����w�
��G�����|M�`veѾmK5��&�І-���>�z�t�:� NM�����|�X�XSqL*��F�g��j�y3�ɷ3@�pĕ=��	�#r��4j��D��oH;a	4�?�ϥ��~a�.2O��'~�$��D6lpJA��?z���s�5����~�Tm���ng�6���f�Ȣ�1]�@U�q2:�&�L$���u&�͖�Q�&¡�T�ٱ�?�ó�+tN�	�������$�H\PW.����9��
����m	�(�A^@	�HE�+��U�񦣤Ĥ���D��2��kb������UVbe8���xq���=L+5\�Gj�E�x���D�s��u�;���e��j���aq���Q���i�t��Y���	]lBH3B��c�,_go��I��қ�eUE�'٤~G@E����
$p��UP��`j�&9?oJ�"	�U�D�&f��h2��>_��Tm�:~T�G�kv.�LA}���!;u�ō�H��������yh�t1�*��CP&ğ6�9:2I�'{���B�u{ͅD�,�� +e��u�L��od �b�Q��)c
����%|y��Uk8+�Z/���/�(�kB�O�"N 4 ��O]��j�:�z�����\)�#7>⋿R���_�Q��T��U,ջp�c���{#ş��+VFk�����U����d�)�u�s�#���"�?F �ū�S>�J�KI4�� ��cflBM����D��_�S�^�St}��*jf��LiT���b��#�fH�llz��b��x(l��W�=���0_�8��3i�-��u2�9����n���q,	D�P'-Dd~��&�����vh:M7��N�I�i�A@��L�~Ã�Q�C�.|��8>�[5s����]�Z�p1��q�t��� (��Lz�ςr��U#��`��9�K(�n|Oа��l�Û�g�z$��g����%}mg��@Is�h�7Q$��r�3wS�m��]�O�{Ѕ��=ǳ#Q���3B�~姉vRq��k�J��@%M���Ċ��&l����:�K|��hL���J_ܛ���&�]Pz��,�Q?��L�r�5ў��c`��$�j~�W]�զ�����٣�*ߦ�����'��ո���Kx�k�9��+#��"�c�s�(�Xn`mtN=��|J_'�٨_,=�����W{��i��_����XW�}]!�J�y�ZJ�hf�x���>ٯJ�E���	=��k�E�؂�s6���D��#�b��.c}�z(���FбĕHF��!X*2Ո'H��50KAU$3���O� Ӊ跷�@�@jv�!�R�ؿ�����Œ�3տc����~�_������>ҾE�iM'g!W�R�=���/��V'RJBf[�d!	\��K����H�ek>\�I���ӫ���J�&=�|��D�d��?8.�&�o6a�)��{�lh<�h��*�b�tq�+�X?}(d/�|�aY��Z�2[�`%Y�:ν"p�p}�x����gGҹ�i�
G��#�C��M���=͑���(5�Q�>��R�4��v�q�%�_+�5.�bv���X���q_�Q�E�2b?)���ʠ�!LyZ���[����	5��f8�?�G33�J,|r45,�[�:?�����d�	���e-:�Ho�k����C��Y�i��l���zu�5��P�	����˿$�^�w�k�FB���yݛ|P��]�Ű� $
����+�^���_�}���5�H
�

Q��g���DyO}=�6VC�}����q����R]�Ï��((��#C` Cv>���U�E��*Uah�m�֞`.0 �+ϓ��L^26�e�����ߣ�j��-���eog1����b�:��q���eΝC�WB�4��rsS5b�&��^�����S��J�S`�����Vl.�[�R���l��Bx����qCRU��>��7���p�q�vG�PW_�R0�yy��C<n��F�!yi��3����8�e0qp�h��f�s�%X����VP��Xf�߹�L=�̚��̒�_Z�v*�F���T�\�l&7�NѶ"'�L�d��96x]���S+X�鑌Y�ĢMuth����	G�[%*���#QG�w�,�sĚ�DWך����}�-9�	Y<u'��f2قzk_�5�W�1߃�#�dCj|�$HBÒp���l�T�	C�-M1Z
m��GV�21���.�x�#滨x�~�c� �=�c�9g��Ц� s��>�UOsȱ�P�RӞ����^��[U��bh)�;!2�â��^\���<i"|���Ed���{<uM7�XC+���O��5���o��7^��^~���T��,�wb�:���;ZV��	&@Qqz�r"��O7��A(㽫B�Ss�&a��Ы��;��wզʻ�b8�m��~���/<��wR���\P���2�
|8�N&d�mh����3��o�@�{߁�5��M���Ҿو����2Uؖxʡb�ջ�vT���Z��Sa>��/��yd�/%�%�n����D����!��z��ݜ9*��ȴ�I;#�Xn*t9eY
W��Hf, ���wE
BǛU�X+k��`�f�兘�Z$M~sN�.���V2�0�ߵe�^w蟀�,(^4�C`?c�� �-�p�6��Q��M����/�]��M�5+�p[0��D��EF$�4~'���W�����kr�ƺu��Yro�x<�b*�1��p�5`�e�h�\�/�Sh�0���.�$FA�`O�M0�([6r��2sO�/ՠ1|"��:�#;?.f�9$Ѧē(�~��ۺ�O�<�o�����|^��T��ҋ��]A�&�|�W���h+��ГɪqB'u��f�mm�N�w�w�Uz�l��&#@�ww0`Q��,
�Ŭ�6^���mJ��m��y-�ѽ?z�4��E�1��H��f#�^l�z���Rg�]Gّ�&T{��&Լ�cüb�خ-�����gj$D���� hl������ý\�`?t�Z���D�;���ƴ"b��G���tT��A��M3��b�i���o�����j4������K��B�T�a&Eh�2�\
���,��8�|�3�\��������m��p
�c
*�z8	m�s}��[�)E�� �(D�S����^�v����.~?}2��t�	��[o�����`w�[�yo�bn �.��R�e}����E���1۶H?B���h/>iN�"(i�yS�l\�
V���l�1�]�󖺼?O��Ym׊��#��Y��XY۵�M�N�-'�Ti;�P��do�Š�
�i��L��[G��56�����B��.-�7(3�$����1��4�����nBL�W�����C4�"6�^}U�=~6�/����	�L���Z;�t7��l���gz$���C��j"��AV�A�ZN�0H%5p=����#?7�c���kp������!��L�5d6t�֪/ڗq��'�~Z���I�������O���'�c�Twy�u���3�C8��P���2\iiwlj�������*'���`>]�ZY଩������]�%�V��c���k3爎l^9
h���4�O�D���A� B�9���k6�Bu���I"�c�PE��4�tu��O|��&0�C��9H�'�i�T�S��p<�P��^����3P��#���!vb�-4��-/?������1�N��m�͞ ��*���{�M���K1w���a��0�W���*m�+��T�aDlb�ɞ���g�`��q�	{sgd~� ��b�U��|Ԡ�_���a�|U1����-kD1�%��a��6&N�C�b��bp9&7����Q��M���]и7�L2�3�}	���e/T�Q\%�*��Ї�2��˭��q����_�����!'�v�]���Fl�T���|�U��u��Tc�0����ީyz���V_Z�ԏ�V૵���*ݕ�9l���L�h�ծic��ń��9�2�a�3��/ ��p�e�"��ښ.�LF��w�ӧ���\)Y�$�X��.�ؼG%6#�P<��X���V/hi>�
XÀ[s2��<���4ʸ�5eW�5�uEn���t�9�C-�u��M�Ae�ܮ�
Oy�X7������&>�Te4�'3�\Pĉ|�G�t�z�ͩc_h���>�^��;E��sT���T�j��黠2Q�m�ҵ[��i�_��}'�j�f(ĈuU�Ђ��1�K��̮� 5}�׳�P�g�7W�#��7|��33�O]kG�cj*�W�ՕN0�#�#��8 ����t\mʄ�ZbN籍�����҆	�v��8�2|E�v+��־.]Ff�Zb؉
���/2)����z���f-�����wg�� ��k�6�BsO���)�.{G_�� C(�aA��)�`c�re���9��G*��K9��]L��:�*�����e��d��'4��e�-b?��C����?�ڀ8ݓ2�?ǭ1�������c����>e�!ʉ�gOW!���^��%�$.8۫�ʚ
�K�����3����)�L��l����$�����JK(�mw��9N��b���l�\i�c�Q:�E�j����(%[ �0����ߟ�7�z�Ӆ�o�\�q�snŭa")�Zp���!�Ѯi~=���I\�t6���ݳ�#=�%���Ss#C2��/D9��,��>>�k�E��/����j�x&�p�����Nf��aLy]���E4�\��+{���j������B;$�)�Z�ᒾ�if���T��� +��0�j=�o��%%��ξ��S���)-ȡ�u�ȇM&��5rj������ΐ�����j�H��oT,8���9��n�r���6L�K5���r�/!�@���E����2-�j��>�C��b�]���]R'���>�W��:�ǳ�j��A�x)Evd�PS>�@�a���3��C��q����R���Z86��W�B~��q-D��"��Dse��Z���7�q��ޏ�T��Jc� �)=	��O��u�#At����#��~���u�'����v�S�J|��7��a�ozm.o5�s5���L����e�;I�_�6�/|�ZONKʮ5����^��=�ɬ��v'"����7捴=:�u3S�1UMa�-���̢v��*��#�����J���<nrS��#�警>վ<����a8X����Y>cj?�(-Uׇ$蓋�8l���0,�Qyc�{; ��T7�)���	2����+'$�G�٨�S�޽2Y��@zj/�5C��+���B�w��S/
��[�uh�i��:��9�K2S�Pe7s�Joa^�h��@�{�����~�]4���2��p1��j�:��΄�U�$ ��U���/.�Gp,kE���cu�z1����Iel�W�����y�U{왔�<
ث��9i����_�3TJ�+eE�}��*�J��i��iT��=p�����Ĉ�&`��@�֗+#�ǥ�*'��G�6�
{C&�#l�[�S��U8�ϐ���"��/�ۅ�=�֔|f�S�~w��7�ٚ��D-�;�si�aq�cv=.�E��y�/{��QO�e����!� 11���h��w��ƚ�Q������wSK��p�?�Fw��L��
���"yj�A�Z���rh���T��\��*&2c��ع����RnF:��%�=B����Q�E"�<��:���Q�J�2�!�[����m�DYf�4��yˎ�
~O7�G�����Sm�� �kX��'���y��n7���O������i�fsu{O�tn {*#G�4LIo��k�G���i?$y4��hT�Sc��єa	w�Ou�y=%=��EX��
�r�ک�5Y�Bb��y�u�@MU��[����vk�#�v9H�}��'H;bmL2���Rc��.�/Ď'�H��&�E�:���x
�,�ȏzo�+���ȃ�m(p��s�P�(mӢ��@�E���\�p�A����"1�¡��|򎹀����E���o/�.țA�n
����8�N
����S�	~홉X���s�<�l�D�gp����]6Z��0�ڋ >N�bԯh*��t+��qb#�R��#�H\µ�խaY��<B��(�~*���������,��j��pk`�aF���83p��A�m�LY�^b���ԦH=v�`��2]�>k��0x@���}�{�u�Ǫ=[�Nyar�	�5�����n�Ց��P��3�ݫ��iƀ�7��q�y�N��:�ٴ�;� 7JaL+���[U������^���C�a��E��G����f"��O�n�I���*qs��L�S|�G��{)=��R�������k�!�����q271:ɁB�vb�k�UP�[�z��� ����g�j~�f&%Ba�3l������	�l���ל�6�y���1�-�����YM����W�����)6i���'q���3�N�?��c'�~b�H�n%�9�r��[e���ƷB�}��|J�b�l�{��S���ܝJ�Ԛ����eǍp�Pn=jWn��-���3�)/�i���B�!��7���]��2�]�]�{I>�q?�p�¯��m�����l�~PD�l1���"L޲z*����d͌��@���M��)Ȱ��{8��$4�c���@kwӷR�?SР7c��z�~S�3]RB��#pxG_�1�M���8=��V�G�g�=P��]���Y��ߌ^$��
�S��Rk^Z=t�wX �0c�(��"Y�]�tA>��hIh=�Ks���g��s����s�ى�G�b(7��ʵO����gIN*ɒ��'��%�P�z�^b��cpy�A-�A�T�V�/�2}��wxu�?⍵�ç�C�nvtoۍl�Ө�7�s����9#��!u�my�*��,����sEd���"B2�s�o���i�������p6i͗�������š	|?�;D��_�� �7�>l	��ʛMH.�T���'IU��S���5
�ުR�%��KU�\�M��sC&u��a!�A�4U�<���y:�%�b�@����ܸ�}��My^�
��&ލ�uj�o�I~�˦�e�Q�k�<ˉ[.�"�i���"��0N�����Ǽ:�cI_�+sV�֥�JkN%�RD{��.8�M�mu�]&�/�!������/L" ���Dܘ.ǣa��J��C����������-���0�&W����9�y�I�v�m�Wԓ��>,%��]�D�.S�y`7���%��Hor���n�E�4���{V��y9Bq���f忯�ɴ��oHQ��$K�,3 v�RE0{hLi9+<≖��*��� ��~�c�z��������!�jQ<(U��O��V�Q\�=�`.��i⤾H����4���9w��i�d$�����O"&��Íb��*�?��_�q� 
�^�Н)���ITd���z��48�z�T*���hN(/��ί Sx�=%g��{zo�/��E���"44aa"���k����\go`<GL
V�a�.�i���^�g�l��` �#�r>�������:U>���bp�?2���hJc�<�R���Y�u����2�+���}�B��d�}tZL��j�i!�ni��Y�;�ۖ�P�	�+{szb����l�:���v�:)v�FI3'�#�D|�bj9I�F�j�H��	N���r#=#�2J��i�0{
h�89~�P̨�VMm%���$�O�7���h�
��Ml�a���E�*-�k��1���{�5���'�,�޼DQ�۾�c��H�3�"�èX�N��'�����&K���/�6��Tu��DƈQa�����`�m�u����9\-%��CO�~zֵ����Q����P�T4Ct���i��������Z��[XB��is����@������p�-���%��z|�r�"���g#9\E��
��1$�|C0=G��� �
K��!_(�Y���9�4J	,F�^7�{��'{V��(���1�;V�	=�^�� `�E�^:�T{Rb��9�lO�g��s��`��\�#J(J�$���L�PdT5����/ei'ॖN��WѨ�%������0xs�#�q@)B��c�qh���s�i[�gh����Y���H<�=?���n6p=�>���g�ˌ;� �f�.I���,4�>,�>��yX�=g�x�w����1��E�UQ��a.|Z���vU�X��׌Aۼ�ϝ�ϙ�^g|S���T���E�!%�%`��̈�\H��!�g�)��w�V���g.68�Ow�����UӒ�"9�Ag������$��I:X�M�e^��Q�ɇ'����OR�P�֙�����@wڰ%�9L[G���;�?��N�˻��f 5�.��d[#x��z@���k`�U�W��
���Y�z��9̈�2��Ϊ���ߡ�y٘�Η��G�`�����w�K@�Z��uh���^�y�:�G�:��.۸�����>^f�:��yG��4�A�Sje�y����+.�4G���a�|$Jҗb�mB	���h�IG����t��Ǘh��h%3o^�����R-,<P����:7��)M!(R�r
Bbd&�^�!y��t��9%�X=�~�bQ�^"/;j4�W��.������|Lx���"<�;D/�^��~ �%`��Ý�$����iC��B�uZ:�F�y���!Y�ȳ�w�ԯ���b��6�w�d���t�`��0�M$�X���@�%Ɐ�~�����*,
��I��o�M�ߜ|��3�:�F��n�`�!��pHz?���	C��%�`;n�F%�u4���7��!�L��z�Rɞq��fLA�y;P��d�g/0U%� ���8��D��	$`���o�>$C���4F�zL��J�H�(�z �U�7_P��B��x�S�1��q?�n�e�[P����j5~�m�O�կ4��Ŏ��`8+Ҟ���9�Xm��k(7Moy��j�sU������� ]�,=!?I}�H<JA~��[H�\�Iɗ�
�G��f+�ä(E�N������IP���;t;���)�z��I���-a���Hb���1�|v�Cژ��an��NB^b�T�#� �sF�E�,�o������4&0�:�w�����e��]�N_�8���� W�6�\��ˍ�[8��b��@�B�Q2��q��Q��{4G��cūvg��eMߌT��K͞�8���Zb��W~)����u?+��|�m*��e�^�<�쯣�:8�O[�]�����E�}?L��RvX$��1���oT� nG Z�^���u�,��%�H�֡����^��$��s�]��=���`C�
w2�?�[�y�g/���P���9>��j�BQ�eY�FZ��M[��Н��S<HaKc#��c�{���?'%�=[������eU���y�F�B��d_zA�q	ɢ�j�)K��.���V���L�',����x����(^=���S(��B��W���
Mq'�x��!w��;jOC��[|��1�ԏ�S�)�$��$���y1,B,l7�redy�*�ݾ%��~7���O-�>�|2�7F�ȳ[Tn���c��dK�#��
+�ȳ�p�l4�J<��wh�J����PQ�9��xS�EI&.�Ū��vV�J�ĸ�d�R��v3�7ղVK\��wg��Jf�ϕwZ��󕨅
�y+g��?��3������J}��t�+a��h1�	ؑ�ܰ�73�����Œ��J�j�>z�O?/��J��د;:s�#/3?�(I���>��L�<�֡�b�x�*N<P1P�)�1
�&Ņ+�'!��w�@нn��ǫ��G��#%��v؟�(��e�/�?v��'!����t�|�7>Il�z�a{��U+�zӃz�X<���ݥ#����(T�6ȣX�*#�)�B����LK��3݅(/�L��o�y��]8?�+�x���⵹E��K툗��C�c���f�tDE�25xY�⠆w�Q'�C2&�
*-�MwF�V�cB���f:`�d��Wu�`}i���&�4^Fh_`���h��fv�?�!*�ҟ_�R]W@�Pjլѻ�G��801ޒ�s��ȶX1ZJ|{u���.��e�����
�TV�����}o���`�ȶ#�'��cu�붞=��Y�?�6��&��>NF���8�]�VC#���X���^e�d��w���AK�����z^]>x$AEiG$=C�@���g�:V_����ya���ڶ�F�v"����*f�'��U�g?��L*{����,v ,G����
v��jPs�AQ�T)g�%fp_8�!�q(Z�eB�ȁO+<(�e��7@�dS��!è驠��u�\8!�.�QP}�hi=U^����	1�M
V��j�A>C�mQ�7�������#1�\5=H`a[�W�w$� ���*V&�VQH%��D�6�
Ͱ�';J��*I$:n iI4��3Q!y��\S�}�' _�N\FY�Ν~�~�����ܗ�;ZiH�<����
�Q�zDK��kEM��~V��7��8���LYr��E�j�KRa�$������e�&/y�<&n��ٱU��1X2G	�$�J1�,�61s3��g�+Զ�,F(Ք�{�J���O��2-�������]�­_n���0�5�$a���G��������X�&��_�4��^���$�ܟ��̎,{~`���|e����j�X[�����ʒ����[<��5�M��������P~�%��x+��PJ����Ȱ�&h?]}������=��N�ڦg�&�R��lپ�>�̪ ����Aq'H)�(n�`��=�'��M�/I���o[�ǅb:�#Ԫ��T�إ|�	��D��z�I[�n�����iJ�	.c�a�o���|�w�~Tg�m��&K�s����#˩�XW�P��TY�M$*c$�l�(tu� ��8��
(_v�#����,l=�*���bΞ�&ᔢ��zL�?�2v�4���d�y���B�iZm�+����'o�+��6���(�GeV�d��CE՘w��k�^����wN�.ù%'��X�i������`^L�3�B_M��2���v���a�م�V��D�~Np�'�<�QH���&�Ri�Q������.��܆���lQP1G��^Ŀ�ܤ+�[��
Y~UX&�V����R��r�3N�/������I��
�_�8����_�yf����㳹� zۦ�����z�1#@���7'pɖ0cV� d]�t9��ݍ'�`����p��\)=���.��E�x�[A;�����c!�#G��Y�m���3�M�(�9z�d+���bK��۫�!/H�"��ԅ�-�ԛq/R�1ip�{��/��D�;�8�.�0؆�v�4�@'t��j�;����
[�7�!m*y���utq�%��׈�p�#W�P0�ʧ���ܙ�U,������8L�?ɋk�p5'��$<fe%��H>Oåbyw Tzww���,iѹl'$�\z�x�]ի��ۘ��=L�䦱K�����}i(BO˙���[���i�R/�!4 ��<��?�o�>���SJ5z�����j�~Ш��Q�����-�Z���Z���4{]���Q�u���+
��5J�e!h�|�w�@���0ʃl�М2/9v��,���{J��$��D�IiR.�*���ڲ����ˍdbkq�?�Qd�����O�<��'����$�Π���߽��]���Ǘ}��k�Rn2>����8@<I2���0����o�VB4�s×|=I?x�����{���O:��Q�3B,��K�(�"�qϻ�y�'��`���$��e\�k�LȏY�p�9:�G�h����M�A�!}wHyo��Y#H���sԮ�"��o��K-����0��}V/PcR���ü㣝����L�r���)xSk�5��Lkw^���p2'�!�z3.y��_E��۠��S���.�����<#R+��[�:#�Hn���UM�6��.Y�Yv�e��"_S�:��D7{�^�6gmk�~#��Q��6-��B.�`[��K���r�_��wa�7*v��7�sS�)NA����YR���Z��0w1.����_r�X��O �T��0|{�#���A�;��ǘ����>y�S�F{�b���1��Ip�����I��Z�ܮ��S}�Ÿ���+|2���Y�e���Uȣ�AA�����S+�4Q���e�w�uX~�#z=��[E�Կk�(��ޭ�.�cc��I�&#ב&%\p���q!�0�Ğߧ�6O�x��e�g���{E�1)ՙ�
n�_��X��P�auE��y��T����\%ol��mE��{��m��e������^�浠d��Ϻ�����jN��gy�/7�^j2F�K4�܈���	�Lk�a�i�'Q�g��kZ.bU�!u��.�Q��*{>_�}�J3&���v{>���9EG�+�M-����t�Zǯ"�J�8�w��{=�N�}���+{���܎�ҸZ�M�B�F�f�5bp��R�K�d~���qo����tus���r��=ZUN��KP� Y�'$���#&�9���'��t� t��@vp`�>h�ۤ�hz
M����=�,H�sH8�Є��=�����n���4H��>�{��HΥ�7�o��¹D\(Z�O�$�G��3����R>��?��!�[{���=�d��S�u��U*��"E�mnx�H��J*}eX�K�{������o�,
j&h��d�-�A�'6�xꎛ�<Z�5����������y�wr�1�?�w�1^j�a&�x<�6�l��B�Z�˔u$����vG�}:>.zY��-��e^X�rx���QL��
@�B��V���q�8\S�.F�!9�/��,mJ�^���V� �U�n&���$i��	I�����_-�g��[۾����4Z<��j�A�:���9I`�x����>]K�|$�:�:*T������Clx`����?N��"ȟ7����2�lz�+�7�^�7��]dy<����Hlҭ�w��,��&f�E,┠KegP�|��� �D���h��O���Z�����h%�WR�Eqx���N�eyWy�Vd;���j�ޓ��Ž�@��2�/ܞ~��}��S�]�"�44]���'�1��f����$��õ��vZ9��&����y�a���LeD�֗ �m�Ly���f��6ͧp��A����<y�Rn�l�	t'�Nܴ�[]�,4Y����$W�yԇ0���r����� T��nx;��I�0Fc�����H�9"�����)�ۏ����O���^�B�m�y�����9ɶ��?<���#i�O.}�������HE���{<�b4��ɕG}3]d�:lՙ��[vW��4H����%S��D@؏����r7�*GZs���s"Q����2�M�W�i%�p`��9<"���s�H�G�G��T���e� ���m�3+�W�|�_���6�_�וd!�7��-�5;��}���l��)s�~#�X ֣�_&��:U�������85pu!�l����Ʃg��^p.�*�2:.��#Il$�����7����G��s�*V}~8�M�̘��Nӯ�t���>�<�<`?z�m���G~77裱s��P:ڀ��أ��C� ���1�`��ۯk 2wNdXpQ6�K��&k�C	M2P��ѭ�8�ҙ�:��o��j
�{���i�'�����J[���S��V^�.
��l��	���8�{�o�� �\de���o�y���gy�
�B�FV�Pq��w�h4$7_�i��c���ϠQ�<v���mO��[x��[[��A}gd��M��_X_z���:���&�-���;7�:4�
��CJ�וpD�4����IY�/ծ�1'W�-��o-l�  �<8BE�6KT[����TH��7�ǔ�R�f��h���N.�P"w�d3Ä��帿�z�\��e{��C��Z'�.ܽD�p|g��y��ο��c�.�7����;��w�����nXEw�K��R��c�x�条�>9�)�'�S0ֵB�$\�(A��1&��=3��x�p8p"�k�z��4�~T��j��k��xR9��m�� .{�L���<H�)�N�G	���i��3h�ư� �Zz�B�Xk�Ni�!�N��j��˴�4y�h��.�i�1�J��bﻐ݋�="�N��N	��V������x
A��M�(Cwa��&�05�ѧ�������U�g�8o
���`��-�v��0�l����x������-�����t�t9�1�}�t��垸��܎��F����S��,�zn���8y��f#�7�	��CR��E�_��t�������1�ĕ�H��0�U$lu��m%4�]8�i��3�i+8kG�c
�=�d]N�'=B-+!*/�?���͎���$����e�LoF3'��4$���ˢC��F�����W�y����&k��Ve��7�_|&�	��~�tw�1`wV�V�^� �c�-��^�R:ѷť�~&U��źE��F)Z���_ ���Sm~s�yw5�b��4���3��<�G�B�|:��1WE�|hN����Z#��*9�IK!����Ŭ�����B7��D1r"�=F�ed��'���Z<����t��'0���V��E�����dk@��J��t6V;AX6�WM�$�R$��O��'1�q5�r�-�c�YOhu+=��?�@������<�G��{N��I�Y5��0+�Ѹ�_#�]s�,�}�;:���
_�w��I1�>�!��%�{̀�o�$��a	��m��i������v���� �	�੤P䶾fu�]�� ��2���zX;W6?I���l����o�cZ30�8N�cٸc]I̪��:����a��gi	}1Q)���a�¡R
�I�'=u0�
��|��X~<���f� c-�h���$��$�N��|N�.��%A�ݚrs&�H�Pk��j��Mg�#B�-�f�Q*L髃��9�W��9�������wZt���uj�9�V��v7Ce`Dґ�o��K*Fͽ\W]���	(��q�Dpg����0�U}��)T��`��X�#r�-�(N؟������9^� ���O(���x�ӑ��q�N.�U�<��#יU_&N����"K)M N�{�[?+K��(���x<9����;���m���3��՝�»\ڪ��i;�(I�>����ؖ�1�0H�)	��6s\{��٘a�;N)c7GSsx#�L
�A�2�i0]����5'�����Uo�DՁ7�Cd������M�<��3S�jҠ��#)G8>D�H��_���M��,F��עwҙ��-k%�L�M`3G�u�ب����	�c�@t�W���6ˆ�k2x�!F����B9G��_R>�L���^�O�TΖ�;e͋�"�����"��R��`@Ї.G��A��	0�ܐ�gė�K�B�}6-�Sf@E,hu1�˿�3^lCo�5+���Q�DE*��7'�H�vl�JVZp�c�{�	�iƢI.����j�Z����S�[��E�hg��y��?��v�m�����'n\�+�c�'DyX���=��%��Q0�Py�_�<��(b��"�]|��%���Y�y�8-��#����%�i�GN4��G"{����z����Ru�h��3��%,0�kg���.�q��u��h�y�>3S ʨ�v��ul�&��j/#��� ���[��.�^��1��0DOڀ�l�5�XzD��"����o��>#�l�hD_
��&����;�6Ů1�>@������&/��y�6H�L`��������'� ffs:5-��d�pXRO�Ȁ[!φm��ʋ�Zh\��.��%��*��0hzb�c�?{��i�Oq�e���2pT߂�"�|���?��"h��aپw�������2D������;�2���Uyd����\����I#\Cs -�ݽ�@j>�|c��=���D�ʖq2]�p'�[�L=�o�C��q���)\l��Nu ��d����S�j+yiY�T#k�&��v�
����!>ȩ<���B�	$.���r���6"��	�γ43��ky���!wؔ�x ����0�5�7�0$!�q��jYRv�t4�� R9}0�آ�mjg����[z���blShh��m��Z�d�_ey6@�	��+yP��� 󮮂�߻vCq
�S]e6F;K�fT��)w^���;-2����*����Ү�t;M�pOՔ�%��`�tMM%Z~�j�ݜ�8[�`������|x��T�p�/x%ϵ6@����s	�AK�%Cq�n��K��>�4d(sd��1Ps��Ks�u_��}|�aۇt[?�P���"�W9��KkN�|#�%�2�}\�~�'�kǾ��D�z�@�*�>�A����1�z���çĖ>O�nL��R<��Ҙ=o\��l��9ct�⭞�g5:z�g���{i����9=�r裐x���\s
�Bp�=�#x��&�c�P:�1�7t�1��3�Cڧs.�n%���D��^;p��quNw�'q����W�`V�~ͱ>��VQUA���Ő��R!�W�W��߆m��|�-�L7�����.�5��ɲ=���t|͵��k,�w�iY�#��1SQ�� 8��nk��Y���;q����뺐������X�;�c���َzt�a��绕A�7@{)}\�5+�v[}���xN�B���bu��݂���[��I�$}�Y��g�%�z}}АG�h�X�ﳳƷL ���9�G6/v6"-���K����1 �=��+��ߔ�W#�T&�w�T��v��J%�N�(!*_����C�l[�"�����۶�:�����s���w�l�����R6�x�v%%�{�r�3qY��t��X�$u�2+��M]�~ƺbg�9� ���}�tj�oD�͕��QN�a�!X���F�~D�^k6���M��*�=I�>7��|�ݏM|��#��+�;/i��&�µ]x:,r9��S�0�˼L?X�'�+����טô�K����b�ɟ9�zu����c��|�Un�#��'��e�h���b�g@8?�"s�	!eՎ�xN�h I�^[�o�������}[Y���-�B�?��BÖu����zM�M@xi7w`(���;��F짆A/,�,e��)��Б�;b����n:���w��Y!�a�.��2��÷�4O�q���Q��Q�W8�k��Dvr�-<g����w~����������[>���߀�zq��������P���B,�蕖�YH��Q�k�U���M��4M�7�a����f!�������f�C/a,ׂ��!�wow���#���%�\�򱸬'/���h:���{t����h��l�og��4��#%�]�ps���{�[q������H$>�|$}�B11l!=�Y���dW�u/�{=������f-Dt��N�5�bM�f� �n��C�&⛯3�_.ܺ
�g�G�Q��>UM��[~��ٝ:�m�&��,���"_���ø2�H$,jҘ�{�j���DR���ȖS�0R��P�IϽ�ぢ�A✿�R��c?x�[��9��l�t�	��*jy/I�i�!��Ycq�k�y;Qc1S��z�p�-B�&���,��jZ'O�s��A����� ѹ�fp�v��y��rtpM�x\Y�mv/*��9�� ���K&�*J�{y`2�rm���
�eȎ���� [	�,S���!$s(�y�� �m�7�>�z���$x��ɭ��ON�{�3������)C�hz]`�	�������h7 p��}îgkL
m2�����~���%>ND���t�=ƃ��H޴�n�x&-ZZ���NM�d�/�)[���Gւ��xXnsz�%M� ����!��0,^7g&����GU�58R�N��L����*�(���[N|��KD^�7k�B5�����T�W��۬ꃦ�fD�@�3�yL���c���Gm�4�U4�ȡ}"�s
���a�%{��7���;�٩�+��zDݱ�E�{s����G�L���s�h�8CG��a���/W���$��2ꊫ:���!sIaF>yL?y���1��k��ߞ��@;l��*�I��]Ϭ���&�"�No+�mk�������gC��1�hN #��$���'�׊�b;L?Q���X�iA:��ۑL[�ߍ�-�t�a5�C
����<��,��Z4���)��Iws�8y<Y�h>��"���tQ{��H�����~K�<(��vs�p�?W`K�G�aʲ{|��|l��4朋]qWK�������cl.m�J��VI1��ˢ���ju�Xw"m�Wl�@��.*ag1,�������������ɏ���F�{�|ম��G��@�ѳo�4�mD򜕶d�j)FJ�sN�O5F_J�g�^�gh����W�޴����L����.�l#�q@]u�\N��'UM�g����ps���;�7�C��Y�N�	�+Q�y�H�0"S�Ԥ��dp/�&���	�V����>{��A!��Y�����
c����f��c�0��J�~l���l0�/�x,,�EW'�Nu���S��LmOW��3�B����0�S����k�����s���e�߷2и<��h�N�C!���K�����bcΛ� �],��B��?�g�A\:Y��T$����I���T��/	�k��A���? x�-����ơH��G�+�N#}ȴ��=X!;��)���ܚ�@D�0<�!���#��i'��c$�}{��M�Y����9�/�9	 �A5Q1��	c�VQpX�U���ԇꂠ�B��Cv\d:@��d�E�  �Q4��7�;+*�����"W��Tm��n�C�JT����]$�b*�� �����vc���\�8g<�^k����{�6	&�AdkR��:���7P��{�X��N�-2��"����H)A�<�����
�R�S�t,l��w�Jg��ϥ�%P�q.`�܏�"������g�����]��ސ��
l������{�z�e4ݕk�S
5�d����'��~o�o��X���_/�ecr��A�'zk�&-�;QH���Q��xݭpS@�+���,�3�1D��PO�Va�����A�[ �.6?�Q	��,yI�x�^�ÒN��nnQ�$�8�;(ӼU|�z9���Z�j�u�?0.F/���L�9�q�����)�+Rj2!���mD
�����[_+�܎>.�o�_��y������ԫ|d���=�%�$��m�f}d}Y�L���a�/�5�yp�}v� �5�ڇ��n����=�@�1
@��nm� �B��h3�Z��1���|DZ��g��v������+��[<%)F%`C��۶<;��fK_�Z>��ڵg��Z��FH䣝�[I��r��n�[�F�K���9�	�zhEI��ζh���&�&�='ڒ����\Gyy ��1.ٞ��;��v��d)y��W1M�:o�
fJ�����q���p�+*R��G.������]Р4��\�~�R>c�����0�i�3�H~���u�-P�҈M���ރhXX[���ro���/M��c�z��3i�D�(%����IUV��u�X�h@�����=/�I����$�N�W���Wix,�}le�K^�%����e���#I��^עuf�Č�ҥq�T�x�"��<K�����O?&���u���"�[#�ܞ��Aۚ6{<{�]�����_k�Iw�X~�m%�E�&������}� A_d!�"�P�i��]Q�]GGj���@�r�6h#���R����k����K�i4?�]#�c'��җbo���,���vc�y�����V�g4�)h��~�!}�ݼ�$Q�(R��2`7\g;Z�-��$�O܎:�!6ypo}E����{m����J�0pt��YN�������Q��|N�^���ؒE���Ԓ�,@���LQ)Z80�r8�U�G���}�#��@�b]�Q���(�"�|P�V�"�~K� ���Ds��|��}b�C�v�=u�̸����#-h�9�{�u���Б�s�ϛ~!U�`��;�h ݅�v	nב��+QA5D�JT��`����F�.2�s�&�p"�ke�*`�A��yw�e���aӗ�Cs�Y"V�Y��G�9\S����M�gӼD-m~�Rmnh����:t�2[�t�D��6����]��/r�ZP�^�يC[���z
��YC��z��*�+��F�f������ �Fa�]A�rO,�R�+�� ���N�-�i����f�ap�E��#d�����f�$��!)�,xc���y�sp�}g��8q�t&�N۹]o�8��̽�3_9��4G��a}b$�
�`��7Jz`��QfZ��`�r�N�q�`�}<E����g�X{�p���Z��l?�Bh�1�L3_�
������g�ȳ+�˛�E
uh����K)oб[A �[�Yf��	*HM��g�}�S�b��h�.J��)�s5"�)�/��r�8u��.�SMQ��_���@��V����yޫx�*�Lb6O�K�֕�;Eb��<��r�_�؇���V�C	�����%��y�8ո�E1��ޜ�,d�<P7f���k�3��8��e��O��	U�v�0]s�t+���C�d�"aK�m1�s�t�.���� �g00a���&�ꀞ�$� H>���,�w���C)������c;���D�O��8@1eu2�U�� ��{lf�"�S@Ve��kXŷc���n]�5e�p�7�F���"p3��։K�v �p�7��}�t�	����݄^s�b��a��a9J*�	��C8��������Hc9�H��ͩ�9)Wmߒ7[���$���	0d?�)U�~�u'�J2���&�/�K0����/�5��Қ�(�Ѷi�϶1����k�' ����T�(�����$�w�D/T}�+��H��pmE���w$�q�/�א��l��#^�Ԕ�e�A�zË.d��3Ob(@��%��aE.[L���Y�D�_ Y7e�o���YQ�A�<SU��������aq������Q����n`O��U>�ڬ��S<[�,G�("��~��$9��.Hy�XP�f��_�])+O����)Y�~�Ve=
�������U3J��Ix����W)e�D?lā5Aj<�aũ�2+ç���g��c���ུ��.F�8|m!�1�_\r0��U�2�^��	�] }-t;��늾��5z,��l�vܬ<^��S07�-�<lM*��/p��`e���xn�]!泴��ڣ��b)ʛg��~�f���g�HPx�����	��K~օ6�q�o�|o�~����̋a�@m��ˊb��RO����E�@f#7Ν}��UJ���oj+��̖��ф]������z��+����6��!�V9��r���^
��8��ݝ18le��%��;:��ڏ����ED6��\���Ξ����W�=����V?���A���H��<�k��7l���jk���.M����8�6�UI[��rҬ,���1�^��̎ynܧ�-�ޗ�ʃ������{u������K1�o����y�9h5����Q�90�~t�����>�{`�P'w=^�ن�1O��E�n{D_�+�Ph����7�j�9��W�9�4�V#=�DzW�#&O�:����T�_�^#��-h�Jɩ�ա�̌�I��Cc��zd�u�heآ^�,�ކ;ۢ1$_�W�{d+n��g���'n�!�(X%.�C$��+;��9n��[�ܨ�n�@�/�?ql���f��l��@A����! k�}�
Z�}׻��^�Y;���d��FӁ��\����d "ub.��I{��ۇj�������;��`���>�\8d(�4S�I��:/����#�t�K�P#��F��� ��!ɷ ��v&�m,aA;�sk�.�m^}o���I���ϭ��F{��Ô�F��Z/���|�۳#��Ǿ�/��,ꨩ�6JדG�v���J�d	��{	�j��/�����3WIy��I�րM$��>�أ��2t��������8��P5���;� e�㏒޻�Zy\����zO�Z?K��ǑY�Hd�9�����k�!|�w�#?�n����^��B�n�o"e-��U�	���!�7i�\(̄K���^�f(3D�X� W�~@GAV�	�H܂8��׶�
��γ%	�"�����51��dD��#��J�:��Z���3JW>�h��7�ǥ�wn����}5�ձ���`���
lb���4�^�w�M�a�i��>�=��5H��E�7����xb\�Ir��ԑ�8�H�y�] TaB >o���c��ac�o:r��\��o�U�wer[7���wbd�j��;X��}P6S�z���nEm��k;�!-o���iT�G%��#��X�,��g�K�]����%ޖ����0؝��X������� ������f���y�;.���tӱ[��u`����� u�^�&_�}KBk���ᴒƳ�^H�.���כ׳�9</�x\,���ݟV&��)��q���tH���iq�A
��9'D�1�Y�a+���:�V�C�L�E�����/RЭ�z֣�' ��N�n���m�ID�8L�y"B[�.)�3B�O_fY(˔X4��T���f�Ƞ��NK�X���4p�)Sđ-��4���R�d��C�dp����,o'	��h�Ӊ�^wƴz�,:��~ysa�����a� F�s�y��h����@�2/Ф���*�k���<^S�ǘ�g��p�*�(�h��WhЧ�3��L)�eY�qK�,��`q�,�u4���+�}^�tk���ݦb�t���D�>ʇXPfk��Tl�p���B��)h�)�
�i����*�IUp��տ��h��8RTo�)��t�Ք@}���)�1*#<��S�� �g��A0#��mm�h��I�B�;��gu�z�:��<A����(.>d�W�{���O�K�ݏ� ���UZ �݄͊+��wF��C�z�x$���D|���T�b��7K�ȉ� ��c"�`�п#�+�U��L�1��v~b��Odo���IɤK4e�?C��j�e1��Ss�\�) �>�S��@g	�3Z���F��\�ف��dB@�Xe�����R*)!f"�����xV���y�%��׶A��37r|�����PP�(��j<��ӃX^��
/X��xP�A�P��C'NLj�T$6�qv3m�J��N��Z���~B�s|JE0����?#,A��J}N��B�n���˅����X��-�g��?�;�'ء��F=P��G3��I���r����X���(���5��K^rt�j��@����+��tH(�����5���;�}R�U9�� Z�:xLl��ˠH�
��
���RÂ ����Zs��v��86��f3���e�3j
��9�)��=U4�|��p,^X��u%�F(-M��.��,=���,����xLk^�T6;�+�t*� ]�˗�͖)�j���		9�%�A"�E�C��Z�(�^IYd�0��� j�l��Ľ�����{�&�Z�x\��p�4K�"�Ip�V�Yl4䤇Z�MQI�[pUP����x;B8M�2s?l$�L;�R�����l��i'����9��8H#�"����VF@ZK%���;���1���k��X���K�'[����.�f�<����z��3�ϣ�qL����}�8f������1�����#]@�2k؁d�[�н���0�7*+��u��dJ����-U��1i�$�)�9��IV��!*����W%�5��@�kMk�C���?��
d����T4Ӛ�|]��歂aEI�2R`��w������Jd�:;L�	��!!d���+ĂA���af*LMcQ%&S��v �CM�_bK˔n����̸��DpX�9É�����q�ɤ*b�΅*pc�����J�T��pz�%�s�X��Jx�u� ��,r�#(;���3Fǃ�y��,6�/���_JO5}ž���?$;fz<�dD�'q��䆗٪Xތ�Ih��$�6W4(��l�o�L�Ut]���nvB��[�>L��c���P0�X��9�.�箇��_k.���Λj�^<|�;������$��.-I͆oBo|�{����H�[�ޮ�3nRn&�}5t���oM�0K�[CS����ʒ�(����&�إ�9i����j�=��z�Sam)�P���}�-�Y8���$N�=�
OO�ݍ��)G���{	s�Xl��bP��ק����8=��^̿���݄S��>l�%�ua�&EH�3m���w�I9��i�~*�҃���Ŕ�˰��j
5�FC�8�8����� �k�X�|v�-(�r�;����7\G`��n�-��|>���1��G�:�_(OU��u��� H���8G��r�p���������m�=�ʒ��b�,�R�w^��ύ<)D���3*y���'6���(xW<7�+@٨�^'"Jʺ/���;A��O;(�q�K.2'�4�;�F1�G�$:ǲ�Y?:z�5&*1s��N� %�p,UH��|�➏�zI�a�豏귟�)��H$�l3�s�1���8�� cJ]y&d�&��Ʊr�T̠�c�8�K|�]Kt+͉��{i]�+A��ڳ��ɶ�����:��V<�d�y8�X��#U�P|� M[ۮP���/B,��8"vu��>TY�YQ�hû��X���FA�XU��>z��V�����m�l��'���Քp����K쩆J������W�T�[����.�%�TN�4���8{+!m���:o���!�Cqǵ*����7��d���`�Z�W��H8~x��
����C��������}B���|���FgkG�KJD"��W�l�����T��	���n2z4�'���~H]��)�o�֐�Z��򱚇��U��b��f�o�τ�9.�J�l��;��1W��
��p_9�ξ���쎉����@3��!���-�{V�%T.����5i�:Qx88=Ɠ$�d+ �)ԝ;5"%�WeA����������	iҵ�j1���a�SPߤ� J�6A������&X����l��u$B'3�+TF�TD�avnc�I�E�{=��Z����:]�~���+�I#��%�7~O�V_*��J*Nӎ��`_����d���Nי� BF_�ne'T\a�w�p�4~�M����p��.]�''��`��h������T�	�:ͽ74eJ�$�2R9V�w>��G����pY
~s<5ԇ�Rt�|����B��
���1G����{�M�t2�aٖ9��~qH\*0C+{�S��C�	��G�ɮ|%��\�p�Y��!qZ�?�Q���!��0Z���N�i���B�]���"~�V<)w�eIE���D�FS�ܰ�/��P�U�,�Y9}FLH�S쩔Xڠ*�`���6�����xF}
�̱�N��p�J�H�sm@��U��A�t�+{|��7���e���/�T`��3�_�@�N������'���r���e�R�ߌݹ��N�~ˬ�3Jj�����<���E�DiQ��H�R���Zn�1�j]���$�}��l{�.�sHNF�L&~ue�!�n�>at��:�7�],w�E�� �g��):!]�(~�����e5�|zZ	��rB�4�X�̼(�
F��q��������; �ޔ��j@���X>�X*�����A&zf1��x�A���gM}�Ԙ�,:}�#E�^{��o���;P�ky�S�ꉆ���w@�@�k�GI���p�q#1��0G�3g7H���/� n�����h�a>�J#�El�@�ݒ���6��G�����qj�Y�k��.iČG#+���'��-�1DcIl����;���
��/�֋�I'�@r�2��>42;���%�� �kKrz���ߖ��icak~q!ϗ���^�D���K��yC��*3�Wkl��j�XWAi�ᤨt�ߊ�u_J�hi�
QԴ	/�5��o��|���_�/f�4�_Ƭ�����g�dm���h{��_)h5��ȿ&64�zb�<�Ҭ3��}'2w�7X���l����$�Tl
4�Iz�z�i�����_'0���Ev�-o����s=+T�C�-���b��r�7���C�d�%1Ѫ��X�9�:{��� ��Y=cbF�{Gg�,����=|�6݄S����``����y�ȗ���o���E�)��a�5aE=d�Z�l���5hRX�4�z�A,-̥T�=NK"oD����`Y�nZԅ$�h��A���L�U�q� ҿg6�B����V_��9�4�
F����x�C̉{AD�4?�Vn�s�~Qk�Zl�[�ܼ�e�ʈ�
��$�����N�u���?б��3$Ǯ�Ug���D�mʜyJ����#$.q��#o"0Y��N}8�f'��kp��M�$�\XBX�yX��R#�:; �<�73d�ܺ
\lC+'!�p��Yo�M`T���]�Q�#��W0au��m,�	A��B:3�EX����~�m�|��,�c��_zh�ҥv���hd^��ޓ�;�?f�:DeW��'l�k�yqn����9�e޻yM�}����h��T���{�o`z ��c?x@-c�A��Q�3J������D���X/���{ð�����i7�g��F#I�0��~�b�|��"J?oYw�<�cM�v;-,^�I�D^�98pN�i����́�!3\�fW:��.��rp��QH~ŉ�)� R����Kz�x﹖�E���:4s�E�_3�%-'fqeU��l	�O������X`Mբ|����̳�!��� v�����tn���
u�$��������bl�s�~�ՔkG��1/B�g����"�`��e�k�:ߥ�q���܋_��4[1�آ�O:��,`H�i	�u��X�rN.��(�1���,W����R(�s|��������OY���[s���~�]����[Q���:�q�6���ry&�%S�I�}Fx�⢈�'-U��T�N�Ըi�vn�6�_�CQJ*��0������M-���V�.fx�OQ^�vN � �Ɩ�"KV\lN(�oż�c"��� ��ñ�*�5��rH�R��B�b�3P�y%|�t!#�ߵ�l��^oʉP����:�B�o�H�]9$���G�,� �H���V��р�a;��BX,�TF�dYyOB�_��9�V�fF�Jz�֏~&�P��(�B��;���Ԍ�r���P��)�����/�\�FQ�~"r�7%��h���iZOگf��w�A�S{YTi��߃V5JT�&%�߾-n����U?_�nuϬ�9�cSt֒9��+)���Ǡ�j��-EnCV�����7k�ITf���ghK��*C hֲ��S�je;��k�����fxR:�)����5,@-WhꞜ�)��491S^���>���:���}����C՞�6�6�T�E|ǹ�˧�7�M=�[q/r��%���,_`���=�VK��a&	~B*y5B�F�:�K�/������;��t�vF�̦�`i�SIP�ly����B�{<���.��<�?��?��)]U�iV̾P>Y�,�fY�<�<�b��E��7ߋ���m29����vxT�	��y�T�gf9�K� ���ӥ?�e7��>��IF���gN��A�-M�oA�o4�痨(��Y�sp��SE��+���Z'�<*��M�fi7��C�"�$`��ُM�0�����@j�~�����s_��7-F�|>6�Ɛ��GD63�=<;}#�姚��=��٢�呅N�֖Hp�,4IB����a��A��ͻ�������r�D�3�e�E�?�s��_M�1N(�˞IV@�?�����Mh�C��'q��O�y����덳���ݜ��(!���֨x����D�%�\�� ?������UR9"Y���u���B	2��H���jP��V�W��;��y���X���΃@}1�wZ]�c����֩ϭ��=/!�r/�Ǥ�aR±��XvR�{��,� � �bY�J�@M
5^�҉�s�7"Ń!k�HP�X8����+F��I�zr�[��P˟��S�T���|�%ҕ'9W����դ�	W���6�;��e�5,J�V��ycB	��G^��VW���	:��=�Y��W�}�ͺ�BkIR���!��>�fÑ�<@'�|�G�Uy"���2G�����wXTkCkX��k�!��4�b	�o3�>���f��Y��
�~n���N�Pn��	��g�C�g��
�aQ��;��)�L҈0P��������d��FM�^)f��hp�Ý�O�F���[��hf��[���H�����i����c�Z2
���A�\9#ȱˎ��b4c� ��Jhu�b�	�W��{���z*�-���Z�gH����YY:.��o�������wX�]�<_�/���ϓ�l�~��׬X�YW.{�B�|�ox�{̠,�ɿu'�9��{��z��-��FV�ST��hP���$S/��B�����_S��VȎS��J��ϻ8���Q��.�������zp�}�\����x��,H^U�{i�ï҅�[����x �H�d��nEE�h';A�VZ���"����I�	�M��%�%��sr-���b7鵆'TI��0��S��u��.��֛�e�с�����.���?+w�M��ka�P���h�g����e�EJl����C�ZY�|9���׵4��z�nu���k��uT	㫊�R,�1�6�����	8_�f}�jk`��	��C*O?Z�}Bݑ�����3;퐃d����{C�aܻO�k�bGY5P�Jt�)H5�w�V�2���@>ڝ�g=���
�^������>r8��)�sk��j-Ǎ9M'�l�+s�,,ԯ��jgK�����W6�'ƙi�J�}�"��^F���*�s��T
���5��Xa��0��\���'�hFݙ��Ѭe�éBM���+�6*x��æ�g��ـS�-!t\�&�����S�1/�z?�Wz����XQ�{��J��y$�pR^	O���2�� ���Qb�z��%��=P�<7�]̰O���K?�)�]�*�~� 5���W̍V9R�����P�Lq���٠�i����,3�1��a��d�a�r�B�#n#��N�|�%���5;��*�s��n�	)/&�P���x��V=V���4R��Sl�q���:��.�����9�Z���I\���J��X�`��J�+]�b��ݳ�߁���E�_�1��k�W�ǴEc�`�@}�|��R1J����e��_δwё���u,31Ϧ�P����l���<-���QLwV���������͇ u�_E�	���PN0���H|
4P?+2tǺ�J�Ê/��sP*8�i�1�	I��A���S�M��warr`3v8HDF�^`*F��`y�k74��V���/2NXaMuk=<�%�����g�lo�7*�t}���cǞ��`��==Z�v�72���Fc�Wa�f��fh��>Ѷ�#��+_"��U��P�-۪�Jb6=}���^ǟ�x���W�� 9�����V_l	T#�_rJkS���p���g5��h���kq3h*�#7:*5Opj��c�Q~��cz���Vޚ.�����=�=+y�W=��k2��%q���p�1�������:fYq�q�I�x/�im�K��������뿼�q�=�sG'6ZЉl��Y�W�iڰ��u�T���w���[�;GZ�]&A��;5"�5eD���J��z��֮d�(��#]:��V�L	J93p���2����B��=0�+u�!ZZkR�v�ln�O}�d��z�H�!Jߔ�<�ʩF�V�ع,�֡S8
�a�}-0�zKq����m��BI���/�x�J$wd7?�&����o�=�ޓ`u"� ��8+�$�&E{�
�<WС�+1o�c��5@�R���\��o�Ǎ�W����C ��ܜ�V��\���s��;<G���]|S����gg3��Į����0՝�5��W�LM6?�
������wS��杞�׶ƾ�&�/�05+�;���j%��ד�_̘&�w:Fi���5�TU����$�� �_;@9ø���Cת���js�㞺�F�Hk������7��!�7@���%EI���}f��6'������w�~H',��.��#������MkY���1��v:j�r:�dZ�Y��� ���Y��3p�,���P���swv�zPa1�ː��B��y�/ȍx=�ғ}{�|���̊g�<`Nb��iU��6�1o�f+��?���Ȃ��[6�x��/��f�S�аOy�-�7�L�	K���n��̎�|9;z+�Ǆ�Yy�cڷ^V�Z�t� �!�w�g���i
�ּ4�����V���hk��˟�b�Y��[T�����x�W��,��`�;���eN��'+�1f�C>���Y�AH�J/ė$��olsm9�
y��0ZEV� Hj!vC�u�/�^@��-�mA�:<�+1���p_����xVǵp���&�I7���{u�Y)�~"�Ѯ�:& A��E�k����7����K`nǕ�:&�߻�G��ܴ��v�!�~l�r�Zo��+�=!X�/h��J^2G�l���=�g����תd]��i��rn%�U7��J$쵞�Db�-h��L����#-��TXS�:�$�׍}V�Y�8��Y�E���{���2����P&�K�#Dung9O�eI��}e��k6�j P���t9�dX1��%�^$P�V;��n}����z�ز���O}�� �"Z�8��vr,����	yd��`=g�����L�*��(�< 1�/J���	>������f�.X.��Ӱ��ԡ�����O�(*�L6�W���Uӧ�NyzZ�ޚOVX�5����L��4����D�5�̧p����&��zv��u�T��00pN.7�jsN�geG�ז�R>��.:{8��L��EX��e������i?�����g��L���!����Ӈ���+�@e�����`�j�pM,<)�������o�"�+L�C��6�X}��k�'�u�����r�({������`dq:e�$pu��_N�v��H�Q��:�|�Q�J�	��ߕ"$H��{�:�7'��:R#�;����w �<����EU�Uز�jd�����У�����	+��P��`�B��忂|�ǡ�*Bp�!5rP��T��l�Uh��$��i��_���9҅@"#D�X�O��h
��Qh��2��9 "����P4�>�a~�釆�):�;�r�}��H�o>�c͋�hW�t몚��嫣��Fm�F�%�x�����Kx��8y2udszOe���F7��W���q�ۘ��������i�X�ʥ�9�F��Hh���9v�Y�\)V��sa����fa*֜ڮeX/��_�S��ъFlT��n�l��'��uuטS��"<�?*#���0�o�G�윴��L�;����55#0�9�_��!`�2��̨�)��^ӎzc�Ͻu8���ጠ�{����x?�A6y�A��5v�?F@�=Ȅ)ꏵ�kX�#Y���nWX��O��g��3�Rs]��ɴ������G�̱"l��>t)������TT$�f�	��Ga!���۵����A0G���Z�f��i�rh���77\I�O0��E(�{.U��hEΚ�|$�1*�3��Ŵ���_�DlZ/������d����@4o�gP�%1{)&�$ƞ 4;���3|���.��P��Lj�J�u��P9%����Y�Ta؝�K���+�~�.�]#���PBd�4�����5X�������Ol����z�r��8I@z����վ	��qVG�>p�D���ݶML�'݈��(=A�eZR�K�h�t�S�xT�O	j��O��<!�1��Z0�H�����ڝU�{�PS+�}�Sj7���ĳ�٭T7�C�����QJ�M����������H/-[�	ξŞ��b�ݣɍ��q���'༇Ѱj��W�M�Q�r�7�ҺΦ�9�ا��f���=�G�a��j�1�&��=����0&!����[!(V�����Bg�9�V�gB#|g��O�&������ϭ�uY���f�
����Bo��Y���kל�/Gc�=ґ���_ET2�Р%#�C0Ж�K��e��oR�Y�H���- �=�l�L� O-_�L�P<�Ŀ��3��JT�Ԁ�[����9�5�P��wQ�q����@QbZ�uI}
m���dsq�Z��<M�e�L���,�赌+���5���ojg�e{�"x�r/6&8R`�T�s���02L�Y�^|m�r��1�J+���Wx�Ma*H��~��5h�mr��l3oc���Th����>���:A���t�7� ��Zc���ˇN�6�z}m�ig��Y�E9��߇���Z��rSf6��z�9Az��NDb%"�RNq��p�H;����ߥs�1�\QLt��уݻY�'�����\�O������q�A��SZ�W��`��T���-��'#P$�Wdmڣw�BQ�UJ��us�C�d�D�C�m��mca:E����UW����T�'*�Ơ'o+�
���R����x��އ�Wp��$mw��J��Sj�b�;Q6��<�}]� �ճ��lA�XDԽ{T�$�(���Ɨ�zE��ss�x���.V�R⑑<w�:�?)O�_�)B	]�a����9��3cn<�!�m��Bu�G�f J�qhBJ]/��s]d`��3j!f�� >�	T�P�:C��#���X$I��t*�f_@����v����L����ga^Uy�k��} o�lT�57(����,�|��Y]Y*��ͥ�N����gѿ��2�+�Sq���m`?��هc�������D�c�YӋ?/�頴�3J�A�|r�?=R߀���X��%�5c��<1SXrCY�1x��h�%!L]��6?�гF	E�н��_���N96c�j��N$v�*�L~f�˴��E�2P�=3����1��P
G��͈�
�N74�i�-���vW���}��o"�xt�9_�|��v��4�=��W�#G���y�59ޯSqS�h�r�$�cB���ߙ�b��O.-+l�i�cЙ�>�n��p�@�	 ���,h��&.{+��J�Q@� �_̽g�89��
TQ�_����(�k�N��U΋���ˉןOJZD���˪`j��e��|]`�n-/����Db�D���c��N������o��L�*��}�&��6/T�p*w����ƓOtm�<v��.�f;RUJ�EE���]o�E�k3�Zv	��i_g�"W�=����N�̹���c1�"��������X�B�o��u0`X�ϓ{����c^�])�o�����t�͇�J����q�1�A��V�o�B����YR��͋�N*���Ȱ�_���l@3�����&��j���2��j�\Yf؋"#.r.Z5{S��Uز=�wr�0�y��{�{������L�ƪ�?zٷ������C�,��\B]"�Q���T����p��U�F������d��m�:�Rnc���N�x�/{'c������1�&*�'T��Y�0M�2�O�|�a�{���ܜ���z��{o�����{c�d��("�(ˎtEu	�ދv
�_�*�0�n�����K��W�N m\��[K�)Jc�I��0M�
�M��|5N޲+�jRL�f�g_Y�˘9���|�sV���CVL�L����$��S%��!�����N�f֜b�`�� �{�Mq��AEʕI1~܄���x��;|*
�O�A�/+��)؛�@9'��󑎘���}h��L[��L�?sI�����_�ݸ�h]�O�W��O�R�A� P��u� ����JL����k��#j*��]������E�taF]������G��čb����(���b�W�q㌻���Pܑ��3���FG����Rj-+�Y2s�
�3�0��T��ӐPjJ�#�y��5<�%8�y���,�;7ڡ�D�[�Z珲S�NFO/������tv�{Ř���1go��-����G�у�6L�//��������޸���l�T�j�+����
���'�<mр�6<�u�2NU|�ak0��@����4�J($��2̧8��I'�m*STU76�;d�e�ͼ�!�+��@5����t7	zY�hEr���V1�`�E:0�UM����x-�w�鹖�/B�v2%tj���Nqy�������t*�x�n���a(����/<�XLtESJ� I����j߹��$�ߗp ��s�ۇh�X��q�U:���m�u�O/;U�M���Q�2b�y}hhY�_�<��ۖ[�:��4Ol.{�b���JJVF�Jx��}�F}7n]����eIۄY����&$p�-
��1��Ԣn Y #%E���;��D_����5�لoT'SF3+��Q�On��
TDr ]a��Ś��B瞴�B�L��Kn��'R}�Ǐz�I��A�o�4u��W���Z�M0��p'/��jX{/���C�Y�a���r��Y��.�(Ε
�G!�>x�z��Q�>	�)�]U��> ��(v�g<Zf�X��+�СF�=�jD27�)t�>d����mEP�Z,74��zFJ��8�ٰC�K�n����]l9)��ty�/Ĭ/�쥻$J&�0Í�x��ב8�J���_.�@-FlЙ�[�|�d�O�T�z7�{b�\�9�͑@
�L�������юsΊOw>�8\nl6��n��Q�_�;�[������e��� �`oL�v�݇-�!	�g%WfN���@�E�h�cdh�e�9��Ra��UjnQ����C�
��@��Aĝ�j�������S�#=m�x@��7�k<�(l��D��J�R��)Zg'߸4[Oe���Qr &�ΠO�vj��ϑ�-��~����I��4^��[L=λt���,�f�V�� 
W���G��J��%�W��' �0d�J����獴i�N�	^걟���sq^�3�'�/1�� �*0�0�)YF��rP�$B>o�A��e��V�[��b�э̇��`���*%o��Zv��.�lɶ��Q��Qn�h��,���ՕO��[���y���c���r �G8����5��u����/���>_Y���d���4���2��ch̒$v�=��?SH�oٚ��}]��w��>}C��r����T�/�P,	��ծ!�8h�!� l��4� ^��q�yB�[�M�2))+?��8��>!��X���m���I����D�/��ݒ��)��9G��̡e�J�p��er�dlo��#��ٰ�cj�P<f��e�b�ku"9a�@���>���4��>b��B�k��_�>�Rˉ�k�k&v�L��,Z�#�`���rou��Y�BY�.���OY�����
�Y�$b�[ S���u� h�1��0�(�DV���y���0i��!�x>���Ck�`/3?��'lO�����`����"ӥ����\l�!�'��#Byc�z��=�Fu�~�1T_��U�D��������e�l��NN�7�:��w�����5����9�������X��Ң���z�g�o���iNIWQ��v�!���2��텊��� ���3TVG'p�E��ç=��"N�5�� ��ݙ�K�C핡 ��tؔ��@l�x�_WmsU���s�_S\��,�.�$�#kX��}N3�k��0J��ʄ�f�Ml����V�B+�c�Hjݐ�����^aC{O�0=
�ҋ���˂�>�DS�:-�p�S`_�*�����Ƈ �`xs��TnH��Y�E��n��T����69dl��!v's��a����$�i~��n�R�E�@��L�*f{����Ҳ����'N�X@�Ksǚ�i�g��MCKl��bLI$�Poza[͔�R:�*xW���4���ڪ߅��g;e�ܾe���Bi�ʊ�*���T�u�5�퇗L݄09��#��اܤ7�ǏR^��p��~�������M�5��%�P��/r���Lk�ĳA"�d�^z?%1�l��2��SUOڿB���+h�s��A��6�DzU8��oG.��$���c"d���p�Yw������$�4,^����8�TO�5��� �Vt���R�P��;�ғت�����XO9�H��L�Q-C(�x�v[��̘$%A�eg�93k��"�>_ċ߰���X<-fWS����ҳ�h����S@�5�
�6�n�5�դ�������dʸ�����b�8���-5��������q+~������Ȥj_��:���\�ltӱ�1���$O����� nK�'{�J^(L�ꇅ	R�	<��%����$f����[k�}���}����W:��4Z�.J�!�@CA�)��������<��k�W�)̧��+����A�[�d}�gQ�x���d�L���h�Q���	���[^��
��0ݐ�I��x��c�W�xe]���.N���5q(����s���}�[�:��l`1�\n ��0N���\y 7���P�c I��T)(���n&~m��–�!{GS&�tt�2���ɂ��j(d��!�C �����$D�\���2�B
pr�h�HM��X��E+���0�V��$����*�#�B���0��W�����:�����N*�g�K�w���x�9'�ŏ����]��]���K��u�Fɐ>}�<O@�Č�V��8}�s}�daC�MM�ymhi���A�m7�����G������\�j.��?`d]��7�8��_�$a,������@������so4~eO���< �ʺ����H����SN���z�~ʱ��y�H3c@�R.�G���+]o���錙��vx�B��Ga���B�)|TGI��O���Z����$U������'��k�����vΣ]�c7�Y�g@*�3��E�FfD< ���o�pB.�8����$@��V��h'w��������F�ۂ�Ldt��g>Xs��L}%������)ǉk�O#��~�NÝ��(u�2��Z�ͥSNqQ1>vح�8�w*�c,��R��4��p�sn�z��+��z�~�f7ޠPʗ���t��M�r-^.+���q�����^��ux���� �� 8/�-4$&��e����!5��d4�� �8��	l�;���Y� yo��2�x"�K�@ā���|�.����&�t�qP�/L[3q�w�|e��ڻsD�<�����rW�Uі����&��v���z�dx�y,V�i��4Ź���{m^H�Fj���|���D''i0�1��=M�_�EqN?P���E�۟���&����;�FS0>���RQݬ�ޮ��X�#��I���>�܆��m�i�y�C?%������+���;'�@[g���q�4�H@�O��K�M�Ev�9$����
�&녽y@#�9�@ 5�"���B��MnCc ��5�2p@���f������P#`��!�ʛ�X0��ss
����*rt�<n�2�L�� kb:�(��Y ���!�v�Gz��W�'�~�. ����0	A�(��F���,%����;��o�� �\m��0w����
_K�-�-��9��_w.K�a�p�lRe3��y�a���g��L���B~q	lƪ3���c�a���DX��#��ňV�><�հ�MJp����ɉ�2�G�*90���v�wA2c������)?�����B0A�͌��(��∎} 1�Co��*�I��+��#�6<��S�	k��j�H⭂Sk=���p��gD��
)Ѫ���T�*o+xN��V:���!2���C^��hT��.U��Q{�n����ǈ�ya�U��Q��n+�g�TN:!�c���:L[97�X�1t�k�"f��0|�b���bݨ��"��V�Y�Q��y�k�ST��TR'F�:���*K㜸Ү*��F�Uȇwcd9�ގ�g.�oJʡ�6#��&䅕P��>@����^}�g��-7*�Pڤw��u���Q+7�^��,N���h������}�7B�A�p�w��a���c��������C����f*��S���W��v���Gw����B�OV�`b��Zt�����.~鰳��x�B&й�;]�}�CCl�6[�b<��VKO�p�K��S����+N��O~R��|H��еl���A���c��������LxR{���%��j|��\�/��uoז/Q��}P7(�0������(�6㏁O�KNJ ��h|	�1LO��M�V�Hrα��3?�V?�*	W�m�m[�ǆܒ�6{j^��M��d<s�1�j��y$�A�La�6[��C��&�c�j 8kp3~�>�@v���@>t���ȹ��G��6P��B2'��mu��T�Z�7�L��'W7���,����U�-��h�~]UN;�N��)^��!�vkf�>^W~) ��)�y=4ꕣ)���k6�h_��ȃYH��#n/F2}t �6�,��f *��2���I���X��N������8l՗��	����W���/!���#��p���~y0��C��"�"`�x���r��ڠ�/F���=ssGqqg�Цw�j���1I�*���ީV��VG+��'��s��F�:��7���/?*�G���i�L�Z�9mb	@�`=����ϑЩ��E��Oo�%��k�j��v&shC[��d"��T��V��rȯv�AsP	*gaX��([*�<�1ʯ�z���@S�8�K�yuB�I�u���4�T�e��dj�7�X�@ۍ�`�5.�PS��������ބ]=��m!�ݦ�_��."�� ����=���ܙ ��tQ�V|�P%7�T����ns,F4��̿j׏q�y��yx����h��
tߎ�Ѥ!�Eµ7�/m|!]'{1/\�ðB�Yt�_�]}|��y��v���52�㞂PPsh��N�s*��:	0�S�,JD.^?��"���*c����Q��?4p��L�)k)�6�X�pl�>K?\Κ����$>�פVj��Sd�ju��ZnX�JL��n4N�7��fuI�D���6d�П�ˏP;�W��;����3�	��m͗�ƶ�߹�r��
�C�(B'8��Tu�~.�e��h�͔jy���ȏ/�F}�zÁ,��cl��B ��:�#���Ҿ%�V'�oJB�����I������9�0Uo�l�O���D�b�;�@(�Q
���f�I�Q�Q<Bp��AP��+~OS�'M���jZV� WG�&ŋ���ʒ�*�<]m��C�s��]{��`
����:O�	��ٸ�������e�2.7+�q2�u�z�8��ϼ��Xbv��P<���q����D�����'\��m�����I�7�]
����o4E�0�;���G�j$�W嬡GKNfB�Q�n�q>��K_�V���Qݥ����j�����a.�����ך�}�a�sA8���W��I��ý5`��M{A��x*��8��L������#t�z�~��r�f�޼��q{x�Q�bW&Śę�/̈�۔��:������o���./]��K�>!�u�^8�bfP1a�\!CL5�G����fpq޺'��wa��w��͖��4������%s��;ǀ����TsE���4uED�	<b��٤�k����XJp�DH9e����[O��5�N�L_+jE$v�}�A�x|�䘘�ͫ�UK>��.C�i�#�~���3�C�Wd���c��!)k/�MZ�_]����We�x!�9�I�����������I�.cf*N��  ��I,�k���o��iN0ܠ�� �A��FF�mU��
fU�1��ɀ�ѿ�2�!��8?(��p)���\�']�� ��,�;�'fދ��끚�����D�����K9s��J�;2lP`IdL�RsF�2�k�SMjF)Q�ܳ�I��1��Fo�Z�3�$_=
�'������T.S��$�����H�����@rK(�V6��,����8�v:��~�˵co��P�@����N���H� ϥ�K�r�<��-�t��m��V	��b~�~�ǜ��P�x�u�V�����i�6�Y�������!q��{yW���n5/���"v���5K�9�H�W�k�V0A��p��|MT"��$�Xu��+���RzW�,:�<<p ��ó��EcL��߭F�b��o�/Dr�mԧ*\����&��ƶE4�>��'@�@^�ѧ�eO�R?�ـs�ZQ��O�6+V}��ʐ��5�ZNtʨ�g,6�]��u��S�No�zjrM��H�J
��Q�R�������r:L1}��d�24�Y�E�~��c5{�I!�J����*Z�VX�-�>O?��˝vٛ��ƕߨ��<iF��/;��fuE�2�l^���A�A�dLys\#�#�i�:������K{w��Kׄw���H삛��p�a~�X*�6^+4�m![)�n�K�𸪛�/st���t
p��b�D�2ufH����*g�(=&�
v:|��E 6��]�����r����X1��|�'�����@�9�M������ҩ��G��g����-�La�Z�����@�0/��)��V�cu���hW���ڤ@g�t�y�����HS��4�O-U;���P?M���ㅻk�� !���'SH��f4��6!���l�ޣ�����m����:� 3ż��Q��A�_V��$� HQ����{��7����k�[&i�*�b��S���)�f�]�0!�m����ň'��.��cǠ(Cё���px}x��W�t�LH��3�z�I���&U-�qvG�ݾ�2�~2��oN��ەϮ5�U_K�3	Cp����TM�I��.���2�sI 
�D#��~��d�x�^ +��|��)�������Cv�0�F� ���Ns�'����?��C�;����m[hm��ҡ�.�Zi�eC	�c�E��	E0�G-�,�#�q�H�<$�p����ge��le�mE�\L s`��x���J��WO��J��?��T��a�M��Vq	��p���$FQ0���v����5�q��r5ؑ��;X43�Q��	@(L��͛�V:�wubS�:�i���^Ŷ�G	tBr���HI�Ң��po�[h�,��q�Yd4��'�x�������n�~��9��	�^_.iၒ�}�6���=�FxL�bB����Q���^�L�$�=��TI;���JE�۳`>��d,S[�V:���l��(G-���'ʃ���M5�qB�e������.h�Wk�O��P�r�$��R*�g�/b�p�@T�-�NhD�u��cӾ�~���T>�d�'��2Z�Y�zcr8mp���"�2��i��D��	`E�E�`����y�xVa��lj��[�/�/�w�� �y���b����5W��%��GI�QK�����_�sz�#�m�4�p<)N~��W��a
��I^�r]�l�Y�3�c.�n�%���Gi�Ɛ8Ls��XjY���.��ZF�2Wy��5I�[�{��[�#�7��ҕ�E��_�ke��!���A8�x]���URi"�}=����� |ӯ��i���O�G"/� WbqRP���m�|R�/��+�F]N,���Q����9��D_�Kpe��\32�l�� ��5�<�U�Ì�:��TX(�O�l~#+����}I2���IL�X�&*��cz- �����@]![�c�{뵳�{�h�l� hʞ��L���m�
���*zL0=�L�$;��r��������vu8��ʔ������*�٧y_�Ƈ{4%�mc��\�_�Lt�3��x�ύ�uT]G�Sw��٨A��Ԑ�!��c;�e8Q ��	��%�ύT�A�����(��I�fK���"_ι�� ">����)_\���\�ᦕP$�&Y����٫ʍ�`� �d8� 1�y����B�I%v�Mv~��ȉf�%E�U�PX�S��\����	�]��Ln��`4��yS� ��(��a�y��b�����&�6�=Ck�5%]�̵���*H|H�Eh�Z�����T�^=�g�0Ɔ���9��b�S�`)�(f��I�����P7�'{��I�׼re��-��_�K�s����|�h�_�E��8��<�����ū�����������|��2�hRߍ���D lW��.r�����c΋5�y^��Ä��P3g����𘚋��(�Cv-ȃ��[�u�{����QG�#�VC�����u��b�k;n ��r�4c󁣬$gQ��Ԡ�~���&��\�uYN�^CKb�ɴ:�%C������9��8Áɞ?����g�?�\q����+YI�������#��VL�Q�ҵp���?��[�,_�턲�DdP�mITg%�':�e��r�2�V����!����*;9~�!L�F�e���	؁燛B¿�Z}}���Q���r����I�밿CC���%�8�8MP� �j~�,����Z|��'�������Hﭮ���.�nʱN܀S��u���K3.��=�ޏK�W��a�0E-"Uk�^�ֆY�B�1�B���k���k����7T��'I���V�L��g��w�"�h�t���9��"�/5	�U���To㴛�r�+�_�M@(��)\� Bមxg�B��!+�C C�Aae�!�:��QWȲ(��)�*�(�]�*l+�uO�G�}���DL:���|��`�W3�z���Ǜ�vǪ�\�ʍ��jC|����o��N����A� ����H�s�k�2�4�-F����EuI5���=�E���c<��%�C��gxc���>h�C���yR�d�2޻�,Pսr5d�U�J�⛢�|V��_�%�f��:�6�vN���8?�y�����?jZ��P�E*3��2I�rSf�D�I�pɪ�L�/(Z12�����c
�Ģ�_�����z�B~�9��d^=u �ЇS��'���b z��f�f�ؠ4����y#��Z���)_B����̏�B�%{���%���5Z�4$&د:͙0����S�xp��ua��@��&��U���
֡��"A��p�ˤ��o��t���nJ,�
��"ɜkQ�C�����8����#Dڥ����,�4L՚�kM&X�TM�r�FV?�N@xT�-`z�_JEpm�Vu��^K�f�i�>�����V�|�g"���q�=^Wx���A.�O��(�&�$��hW~����M�"9�y�(+E��$��XI�!cFI���K����o�~�,�o�}T�/͢X��ك�"�7����� ��Ѽk����B�U6Ő�JY����`ZC�sX� \�=��[/��7�ϫ�쐖3v�,�ű��#N(�Lp,����'�`�)���[�F����>�Ȧ�G��J��(P��#9!��v�bSBr�G��()�
&���w�d�"��/�cX�d��Q� ��"w+���ib
��.&6� ��mS5бH��O,q�#$v,{W�g�V��&�����B���G�����IU@�CZ
- z�;��X���R������ҿ�D<lN<�e���Jr=�O;��4tUb�� Bm�S7u)6����Up"/ ���G���Jo��to[�l��]>�Ll?	,����+� �".�Ed
�����k�ጷ��|�Ȼ4KY��?S�X�}I7M�q���ZT��[Z��������M�#�~��%$�T_���̫�l�0�"����d"�Ϛ�^��
.���yU�2ϐ�3�Pq���z���W{�.ђ�tk��M%۱����EO1̚��n�h!ˀf�ݳN��nT&�h0A��\��[�ɚK�ڌ�ܪ�sj� <��x��`����6�kK�-��BH�?ec*�71���b�����xh]��ʌ�n1ܓ�3��������p.��z� �4���ܝ�8��I�²�Uu;ߩ~���:��(dk �ң ���c<��ٷ�����6(���!E�t�/�oOEb�+�r�+Ak����N����A@��jC�(��\ϊmKQk�)o��@��-2�Y��a(Q�A�6�텨qoqM/r��5��Xa,�č��Ȓ�e�;�JNΣLR�s���*���m��6g�E��#�����z_2w8բ���Z6�DgX?��@��p88υwsꇔ&�4��.U7�2��N�r�x�XI� �V[�����1�:�
4�K ��� �������咝*A<�D�I��KW<=] �m��(����<�7e���U��p>��I���#��_�����UB��;*-2>9��d�;޳mY�hQ������C�}?���_C��?����d ,x$�Oö� R�%�9����:+q����R�Å����#�1I����Zy~��f��,��Fx�����2v��U�]�!<Q$ŏ� IW�6z�Dr)���R>^���87Ye�u�щ�?���pA�d^����`�md�g����sݑ���x��;0��!��\
�5
>� ^���$�ӯB~RN�ְ_h�I�,����]�`���c�Aj��{]���Ń�'�� I�������IN���V�3�7����8H��m�nldxԸ��(z�8�l����`3���d�$H�bՉƴ	�'�&�_�i�EUoS������h|�D�'�����Lլ�B�}	,S��1#��;�wN��!8��3ٽ8�����PwU�R{d��/���ri0nbq��e3���z8�5E�{�L͓M|�f}�^-���ދ����g�?:�����_)�J����0g�y��!:��t��;��g����BH� ��i�%]꼀v��L=a��$4��&@2F�S`�aP��.{~:}�;D���}m=�O�ie�-#�=M;�/���s�"��y�l�ڑ�I�F2HV���wry�	C���N��i�׼�3�f�� q�O۔�?�p�#i�ֵ���?�t��{�,û_UYY�6�u�L�Ǉ>�GL�﫷Z������B����ac�c�i Xݰ��F��昬�o��˹xsy=~j^LŸ*�g�|ifϰ�.�߯Ù"|h#Hr�`p���6���0��lĺŝikU��@F��I2�PG7T���z��� ��~�d���mNa�#���}(����E-e6�D%a��bvA�b<������&D�+>5�`i�I��ռbH$>�`�`�)�{��c�#�G��9T*��N�>�H+O01�i�S�I����Kxe�{@��uۃq�7���8n���%<��lK��E��r:��z5Mʆ/L��g�� �} ɴ�]�a�K��~$iȢ���B�"�)��' �	��I6����`.Vw��*ʔ@l�)�qVŧ����YDb�S*��@睊�̲��YP�.�a�b�l$nwCR�J�[���D���.Q쳼��"/}{\�Il7�zC��Ty+�3��P�K5�D9|A�Ol��GN�ɶ�����#�� �Ņ�:��'<����WLњ;֋���k$�K����ז�U����� 6GL��A1-�4�N{XL����ln\Sb�%ԮdtP���l�%[k8�ݛ{�+l�#B�.�\~�V<�!8B˭Iq���Y��^��m�pi��7H栔0M�2`|*.$�# �*�֏γ��I���r�Z�ޓOz�]Wc���V>`�I D�9H���Ԋ���j����q���R�Ad�:S�B��9_�O�*��N�#�_�$�D �/D�^)j�¾�p��a�5��������hD��ɗWJ��� E.ĩq_љ�9)�o rŦ-���z4jW�K��E;u�<�w�Ĕ�}�!�o��+#g�����Q�)0�`�����r�פ+M���><�s�4Ɓ5SC���ī <z�m҃�����2Ǭ�R<�*`q����G�/)��g:�>O��7���E�[_2��)���@z[�����w�F�I�/$~�쇵[m���
��4#��'�T�~�Z�#b��j�1Ƨ�_7��	�4�7�He����@�z��<<X�	[fc���\�"M�����Q�:j�� _��}\ܿQs�6r���d_Ӽ����g����!����7�t��Eg ܙ#&E<Ú����>9եQ0�K�uyF_�I������1�XY�}ah�[��dr#���*	$>��H�lΚ�m�P�{��n�����0��d��
��j!J���o����-��;H�����H�}�/m
���Ǝgz�t�J-���ɚ�a���˕��&e���^<5U���n�Ȥe!�̓d �!��\q�$� �2��r�� ڃf�k9	�J��Kg3h���!�tag��5��$�st�bߺ{�*�;�~3Vl�;�7�&�N�iWs��Ns���]�Li<Q�ͅ!��c��	/���@ȟ6�:G'���g�N.�2�������k���60M}l_�;�/��~�i�q�	&n���Ǖ��j6_ߦ�AR&���Y�'��i�W$] ���{�0
�Y�7��Ӻ��Q�P|CIS�V*ɯQ��('9�阬z�,E���&�n����M9� �ػ?Np
��
@�K��	���a�l�0��Y��ZR�9�if�����~�F�v}L,�QW�w��ǼAǄ"`J��`���/	{�m�;��'�`����=
�+םё뵲B_��L���H�z�ɕI� �ՒO�4�[i ��[�p�5�"�r�f�V�D#�Qs��:��0|<?W�!hg�9����DFxXF�����ͦ��ȅ2o��f�#Z���>ľ���L]���� �|a��"�8��V�e���480��^M��߫4�Akr�mr���]�k�S��W=!N�+<4�� wr���
`8���@9���b���3\hy4�*�k=	�£z��������K��T���L�X�{O�Jv�r�Zf��qc�У`T��s%9q����%��,�O���|Q�>�."��XE����櫜!���~6uu�n����3�x�L��@��(w�m� q�j�Ȉ�.���j��6<	�����A�U����HK���7���TՏf��o+,0E�6|������aS��zre?f�XL� MI�����{6�9`�F�-n�"dW����Gpr���9`�034$�E# ��as"$ypf-w�x�s|=�� :��g��ؚ����&�&�u�C,�������ظ��JC��|T���*vW�k�7���\.���X�EF��%L;��;�w�t��P�j���msd����r��a���Z;�i`+�0�~r�Р�;_!���"P�hnؔ���r���e��0������	���~��Q�-|�Nw׵�G=;�{�_��0��o��@:�t(�| �ǯ�a3�h�j3��4T�{��*>�f�&VP�>�b��&���"�}o@�	�o��2���$�����"{��
���恗�7�ݬ:���^��e�EX�s��3����_V���c-k�	I�����6q�ў.M~��©�8�#A6���sƱ�R��'��u}��~�ҁx�J4����RT`��v|7R7!Z�����v�:w��h���1O��i��A�+�E��hm\�Bl�@��_ҸYt��Z�`M^��S�AQ-Z��P�G��[��E�M'��I�0���WV.���]�$�*&�C"��0���V�N�
��4Q��Q9�&֛Q���Mz��VեX��-@�jB�X����m�#�,� �av�~�`�J�iD��X�ӴY����~�����Cf���x@qC�EŢ�1��t����l7"�.��~�-����$E�,�R�lJv���~�f`���eWέe3F�zi��-MQ�fw� �x�(&�I�1_��%�c\K�a�Sܻ>K�m0�o�k�=����cqiv��ˮ��ٚJ�Q�Y�k���4"���:��"A�L�]�o��:<o�Pq�C�Z�w%&^2d����*X�,�s7`m�!q�~DD�*��n�*6HT��Q�߅6�*���]��^T�XL#�B7r��a�<�L�!O��>��i/Jθ�|5Qj�]��&�Qj]\=� ͣ��P���Rme�=�sUo�_O'c)����{b;Da.��_��7_T']b���f�V��B�"^�oW�Ѫ��:�8�s��ş��~��N*��!N��/�^�e��v��T�"�wZC i
T	���ܪ$�H�g'����8���a}��(-8È�m��"�j��F��>IѢ`�������;����a�&��zk"	�����Ja���
�F���Sb��_�(��9����� X�.u�[�P*IN+��֬O�.��dY$���� �l�?Ǚ�kʣ�+��sA|���5c6<���,�ZM�Pw���ï���&C�io�t*ϞJ�T>��}��kV�Ԓ�l�@zK_�?��&K��FcSR��c2���S���ha/�,�!{�[���|��D`�`�Ú�_W-����%��J�A-�O� w0�����^�6%���C��ߏ��y�8�?��ъ3�çcpfW(�k��AV{��P��w5Ņ��q�/���
��Ͱ
]�����HRF�Ł\̒����s"��1m���Ч� �J������K2������^	d���N�Fa� �uZ4K��;��c�ܳ��2^u��v�N�J���ӝ ��X��
�5Q^^1yk�<�F؜\g}�5䞒 g�����^*�Q�
$�6��� �c�jf�?��io�SU�ShN�E{Ǩ����S2�@������T�� ��?�w�$R^|-���Xc���B�uM':��:KP��b�6A���q��kg5�3}�g���s.T�7F�����Ur�(TW&sz�pc)�����Y;�u~$�K�J��y��6M�G�Q
�'�}ޢ�Nt��x������� �֓P�:	^V��oU�p�)cNM�������@��Q"P���� �8G�i��I��J+~�/�~��K��>��@���V�o��#�8�Ggua="{��3�2�|�ڴk�ȂB�~��w:\6���bFK��,����:��H/{p�-l��T�u�m��\��P�~�x�U�� ���2�b���W<ЯVB�H������ӑ*'�΀)��i�Z@��pҏ9f6他fS���d�%�����f/ɰ�5o���p�zW����-bO���A$P����]oʕ?����k.ƕy[�e�'�?�ګl�"ֽ��<�!�����R�ʢŽ��B:�[)5+W��D�RhΠ��<[Jc��/@����n0b�#u�un&0j���7E6�X�(M�}�ݸ�#�҉��k���
A���>"�E{ �1�hHL�%vN?wĦј����A�r K"�oP��ؒ/B��$������V����������r;l�nQ���^.��	M�O���	�1���&<��ı�I��Q�!��g}:�e���� �V;��'�7�EƲ���|c$ҩ���=��؄Ȑ�sх8~B(]�.p�W��M=�x�_��I�����ո�^�}��(ք��Z�8h��2��e�}�r��Ҹby \pX<rRI���W�EP����&|suR��B\�ꌌA��]�9��?�-X���*UR]�l[x�Jۀt��s�Kp!RZ��
"��"��������3�^f��7޲��*j׺��H(�����+h����W�0ڬ|Ӟ��j0s����þBB����� �,?���ǫ-���=]�xw�Qu�x������bLڃ��R������C�^���D0�o�ͳǰ���K��)�~�yW�P�Zf�)�1V�
�ɣ������"$�bo~�)(4��Ǧ�Ӆ��T���/��������**���EY��zQ5�6��sD���0����Usv���S���Wt��f�������f��8�߄&�dѮ%�	����IG������}�w+�E�O�aѣ�z�j��s�e*��}��|���M�$ݡ���ȹtȟݤ��j����3�b���0r���~�ƥ�laR���5w3i,5h��E��zi�#��Z�$%�oo��{ȡh#}z���.��i���i�~-��*�h��v�i�.Ķr�8�4������Bj������].
�L�4;��Gq*��=E�'Hۼo2a$��:2�Ǯ0T�-v+�h�����C����ড়F�.u��ah�_�Q3?��dδ-�������2M��$,I�)�1K�w)�\u�K���`H��H�H�`ɗ����\S�L�/6����ts�ߏY�H�'z��<��M��'���$�2
j-uϦG5�!�Z����zy&�G�Xa���9H
�**(qd���舊���p�I�6"����>.+�?y�9u@h/��큛I}��7L������u1�n��=G��j�Zg+4>A�T��P�����w�!�$*�1?A]l��v
g���| v�uF�in/� �,-ʭ잶�z�H-̏�Jf�~�����h�����������XG"�;����1��~^�f9�����(_�>�&}_��KE����;!��m_���F�
�I��ŵgyz�T��� G�+����x(�&=�c.�8a.�LWe�O�
���'�����C��s��v�$��:�:�q�O�k�9x�KA��]6��Fy�)��rÊ�IQ�'c���,`�O#ʸtՒb,�ɍ�����#[��:(<�I(=�|�I,b�,)�-t����-���ݦ02G����-e"��n�߁J��Hț��wё-%)�x4��Op�/|���b}|�P�}3o=2R��H,? �g��2n4��rx
����Y���U7i;P�JZ�@��TK��[��=��t]ÐLBs]�G[�������WK�9����ba�L"��΃�P� ���L$H��jᮕ�t��l%�A��fߦ�dD�wਆlR�)�<<�+�@I�d|��j~90|)�"?���W@t���.�{P��'�MBڧ�9���(�ګ]Y���;G�;��a�139�㞥�����E�+��q����-@��P0%�R���!J��
�Jb�?
,����'p4O���f�����ßei��B�q�ʻ��P�n-U�.�� t21��(�x[=|Ѐ1+?.Ѱ�j��76M]RW��k{���v�9�)��NC�e���s*��l:`7�Őar�p=�a$a�J�cQ�g�A^8�Ur������X�1�qw�� ��a=�C���]��¿��L�T�ص3A�p@PG%����$�r=
�(S��i�,Z�c�1��%댆��h�T���Ӎ�����u�
'�,�D������C_$i+���
��������/��FPi����q4bؙ;ig��v�9�ܨ�H���F�M�����F˷�Q�0넔8��T \��x�y0O�r ev���g��V|�W%�YƏ��H=e��sh/��:�L�q��K�3��ڠ�+�;[o1�|Oc����-�F�w�:�[\b�����������;%(��A瘧�nQЭx׺�x��rҭA��|Ml�p�ʻ^q.,�V���0����岆�Rs��n�/��qҗ�c��h ����+�s8�'�!��/q4���H�͟�W�?F׽�IOW�z[$�	���Ȉu`�\jV@ 2��y2���iԋL��\(����\;"R
OLx`�8I3&p�\ґ:`��&?�R��}�AQ)\����5PII�(G�����µ.ca�r�6�(��i�K�W\"��]��CA��͓��$�~�����N�?�rLS3��C� gl����Pp�K��s�sHl���& v��-}=w�h��j(��(N�GKP��2}\���Wu ���r]�')�f�V�.����t�n�5����f�K;[ѳT��?���*�Ae�7�kU��D+�pqx��A��m�����ud,��+����c�V�ډW3�>^5��>�㼐�0[��P��u���dqx*Ϝm�����M�
��)�9����	�a���;IUw����
R�?��!i���ߒ�84���?�q�ފ.�K*����ȃ(��|�q�g����������wC�@��ii�&�!{?0�� "u�if��<k��>�+h/ؒ�:`|O�B��s!�+���9�C����ۅu��,*\M ��|�9.�#�)\Rz�"m�����Z4�|G�NF� <V�@#���=���݊��]�@�~�}�6��O%x����|rIArH���|{��ճL�G��Uw��z$��o��
R���\39���;~�Kj>�T�C�T�:����<���ԃ�
��u��pk������ak7�g�6��qR⿢r+P��2��*�  �B�f`���>4��I��6k�휘g��o�݈���JC��;�{��A1x)�bw�ɞE�?m�Ƕ��9)�f~���k%�I�9�P	�4��A������z��m����A��.�?ZuEap��6b�r�9�����	0�
����t��$pS#�����Mη%�:��Ky���98�L��h���y��|7�G��c��W셭R����%В F�;���8�@,2u[��T�e*W�W��y�S'كCP����h�5w�
��ÔYk�& �z�����r��-�k�u^��L/=��Rd�E7��e��M���	�h��|yʣ;R��)�:�r�)����X�Ͱ�}�L�*Apf�O3ŝ�s|N�H>~:+�^!���+n����g�Lv�)����f8�M���
��_�_���4CҊ��C�c�ߕ�&��E �� v��p�{#�ϴ�`�E�:V�v�����p�>�d��Y�?.${�=�d�{�Eּ��VÒ��l�m� ��祤Ҷ^��u����$��W�6��bFܻSMB�ͧ8�U�|���D<�s�
6TU��:�n�lz:�7jK�˥Q��qX����8u�����dO#Z�*"���>�Ù�`X��#�U�K_!�%	���P3寝� �^6A�fݕ��Y�K4s���󓓀°+¯q#��@m��G�h�"�6��ŪNc)�ڏ���������B���ȝ��,C�'ώ�s=�oK?�m~"�X;W߃��v>��)��S1֑4FV�s�|�i��I7^+�Ƿk`F;�>���t��;�LM���p���p��T�킧��2��K9� ��Ӏ�!��]\��W?�\Hm�Ō=Q�a-����\����A�����ݥ*V��N�j��U�ܘ�]]�M0����nW����8CX�MP��
��KV��&����������A��p�oEu��9�$�Q͊1WQ~�E�N��Z�9��x𓵫H�d��u=�����b���*r��ݏδ\mE�]
�Y9x�6����&����[B/#;����nf�3��Z���λn�3��h����b������ �Oz�X�Y�`)��E��G4�ȼ��
��2p��~wПfF��a�̲nʷ@�5_��`D?��ۣ;/K�%,:�7 f����6Ftf�S�)������FV������c�'h��#	Ն�f�%������:tR�f?#��v������i>*n���J��'�gV6�/�i�-C#V!	�M:3�E� �Tq��5-=�\�;D�@�%-Z�� wW��̐��|���Ն��>��=Cw�r�贲 ��=	,
ߡ6V¦��e��}�����뽭^��c.�9�s;��u�D�A�k��lU*�NdxC�<U��=�(�UT�MF��!�\�����+����}q�#��n4����'��'�����[��Z�f��̷���n��e����5Jp��[G�\��W�Q����V��ѻΨp�|�t�K`�n���i{q�WP��|Ab�n	�����E��a@��ҫ8��$�i��<���c/��v��-�vV*��[���8�:	���)���}Z�fJ�]��0f��S�Y����tW�{#ٙ�8���$~�v�~���i��t�ղ�����!���/؉��s� �(?�̄k,�,���Y�
`Th%��FKFR
��%F]W�<�nU�l�I�
2z���=�ė?k�=�8���ͥd/rd��m����G�}����������z���������N�'��r�����O$��-�>l�hD*i����U�����L������n{��فC�����~c��%)�Z+�����r<p���F�g�gV��/������n�Nelrw`�`��X�ď�*���zR�ؠN�9��_zc�>��HxGm;N���p5�����;��aq�q�%�� �5���>���OM�	D�~­ $yFϏ���.|kA�<Jf$�v�3rPU`%��ދ+����w�8�p!.E�� /�h0�ʎ�<6�#%�֢וt��0��Pn0 7���ŸЬ�������4��~�N�S*�`5�Ln���H X�S��)�Z9L��P��_փj+۠37m��H�rv��&ۻ�GM���_�+v&�S���ǳ[Q���*�����;�9����
��%��A���.��O̗�]��<�&��o��8�z��f:��fL��1f�0R��3���=��5}�T��(w��!�x2iE䓾�QO��Ғ:</�7���s��|��PՏ�Al�C/,\�Pg�>	f�0j��N�aO���o_�mT@ꦊ�TnPň,�_���x

�;*�X
:�\���ܶ����OI��aY�~4���J]�}H�c�>�Vee}/��vኈ�ͥ��L��Y+���B��QG�)#�r���'���=؞L;�{C� g��	9�׺v�
Պ����>YoPwj0mؒ�b<�4:���Ȱ�n��i� ۥÆՐ3��?��w��E�r7ףm�62���M�Ȣ6�ٜ��W���F�%�4�7����~
jFd�rL�CS���z쁤�p��d�#�:r{���Wi a�4�D����s�Z�:�j!o!�(���О�lc%I�Ɖ["Bn��-���a�<�x����K�p�7��n��~/t��^����)��o�ѣ��Kn�rN��f�d���.��$�����ϒkY�H�F���f������=٧B��ge�#OYz-s���LjL���Q�+��v��-�g�  �t��o����n���G����^�v���m��������:�w�~MR&��<�yX�$=�=}-�m���������ft��\Kط��WGgl�6��@C*&�������UGD�z6��z�?������H�F��v2Lm�Χ콳[ר~�*�3�$F�D�waYTe�{���[���c(����L��������e�2~�1$p%�I��U�1�ruiXY6�ݐkԒ�5�*�_rB��_��h�"_]?#&�� �86[l�p�@�7/�|�����n������Xa����2�Ǘ:W��6	� aV�v��U��ze�E�cQX�7�R�����'I����v4��<R��vCLJ�E���՛(��B�����ʉ�z΋Jo٨�G��|��ڎEĊ�	0l�����^�?�+��v��bOU��E�H'���xe�|_���������64o�%,����\~��B���e� ��l�ͪR7��Ư�I�Hq�c��I�����e*�nå@}�� ���s���)}��x�ŏ�����ʥQy_?=���,{���O��@��p)#��p����9l���_�)�P��ؽKI�a�̓N<m�N�n���X�q��H���xp|G���+NI�^)���2�pI����HQ����@�N�@����^�6����^�V��}R/z]0��nj��g�m�"ul�1�4�2�;������S�Z����@�������S"j��ό`�Y�%ù��g%K����Mv��K*ş�ڽ��d�z��j�L�4��5#Mw5]W%~4�h�B^O���z(�_��0�Je��6�{{�K<ώ����S��F��F��;�|ॉ�\m~6ϱ2����9�ʗ���A{����ċ�DbD�X�G���VGN�y4��y�.�:˞2�r���m��ߎ�e'�2�x��iJz<U2}�4"X�6#��X�b,CឝDp���"LN�'y���^ȭ4��Sh9��)mU�}K!����Sm��,���	*�� �U�� �ٴ;���t�Z�r�W�i�˩J٢��N*͊y���j�J~dD�n�S>�&��VbX��M�Q�d\��M7��{K:�U���������>,���I��eK^����_%g���t]��<k�-�։*�^]o���+���C���(�9��p��Wg��,`(@@8w䇶��w=1�{urk^��&ǀ�(@�#1~i��py��;.�8�?'��"ɓ�g�錘z}43F�Qʉ�z���,;6A�����{9��vEh��4Ͼ�m��%���t
�ZK���HmI'i1�ZP���<�#w7�1�*�F6���h׶�8��ǲ��b\U�Jd�G�QK��+z�~/ݔ���Y$U���	�d> ���ex*�}�7���шO�jԆ�V/��l�s5�F�(���RT��:��� ���� ��ŶV=�*�A^	YU]x�,Pm0.C��R�ub�9��RyT͹��{����V�ZKe�$l/��)���
�_I��{ŮT����v�6��/x�e
��(ꙭ�3�89,��s���Q�b`�d����M�ˢ�J�I�*�������s�ߒ4L�o/��8_$	���~��q�.->q+�}ܪ�
%k*d�$��R��4A�yOTFNf�m�q+�$��/�g���]7E����S���e�x?^[ȵ�-���� B(.�G�ԍ�Zp�u(�.�LO;n�=�D��5	=x��X�9㑯-@*j҅�#�cFk/��>�Zo�6�N�q��Z\`>����Ϯd�V��ގ�3}��yK���4
G��f
ȯ�|��eƹ�yV:��[�R����޹>��������?�Ru�d�!(uR�AS����w� w��w|�ȪΌe�y9w�1�����Ú-FpY����n�!p��e��YgB���_������E���.\]w���(�����"ֲ"�u�ecAW�%U[�m�5�n�g���휺�B�L���bL��-h"	������U�[<p�����w��Kgb������jU�\�a���e� P� O�W��J��`]�ؑ\T�'mב{��G��8��Msq>e��p\`Hv<)��2����0{�PN��*�48~_�+����zYҝ��N@�9D�uW<�}]*�J��g��L�^�λ���īx���i�~ħ猳#O����/��:�3����4?L���z�ۡ�}�?# ڄ�?��T�x���v>ݳ�P�a�l)�/��Y����CS�e-��au�W�c�]5&��Z�~�
�	f��`6��s��bU�ԇ|�XA2�[+�z����Jc{k�غ9>�ů:۫����b�Ilm�78�i`B�O��MG'�[J3('�$�w�0n��舋x�����E�T�U����6]�E@��|�}��j�M���g�U��c!g:ե�
�����`;B�[�Ba�5�3lߖ5[��sX����n�鿸�t���J����(�i��Nw�HI�3!�������TR?�2B�f�K(-�q�OUX��&
�gX�G�D6cwe|�W��I"��f GOyb=�槞�9FKS��\��R�ƥ�>��q�4�m5g6S2���YR�y
1�U*�+D|1n�0�Pop>qT��5dF����� ��Ӿc��!a�9�輍{խ2�2�r,�j�A�!�k_?i�<Y|�"�q�l��{��I�FH9)�$�Q�-}�6�j�� -�C�n�k��ąù�剗e��*n�4W�c�i+���L<�|у^�<������=��5�Ĉ�|q����	��}ĨG�Ϡ�"\#�v���Ȥ�����/�ȡ_�%a��oX�tch��"��h���z4�v(gn
ub��'Y%K����9�#���p�������f�ڄ0����L�
��OD�D� �.M�ۭ�&��hl-���;ĭn�k�!($����4ۗ$mcf�4f��n�ϱ�������}��?ї?Y[��t�z���ІLs�jN$$�Ȅ�O#�9�32������щ��w���"���͋�� �!Zt;��,G�B�f?<�5���9�;���!d輛v~��nց(�'�<n5�&�y�j�c]�10�'���U�*z@n�j�f)��gͪܯ�N��8r�åL$>J�b�f���q�@U`�c6*��~z��#X�Z�@�҆��S�iL�ߥ)�ccab^|9i��E3�K�Kh�����5~��!9���d.?�%G4�V~��k*�Q�i��E�0�s��o�;�� J����ؙ�r�U���F\�;�k���m�TM ^`Tv�F(w�?�z��
|�f�B��GDl��A'��Lud�Ia�9����91��FG�C��9*.�d>2s�s���	�����$"�*��P#D�L��b�(3Eܿ�q�=�H<r�!t��6J�}v��
_�'���~�Ui7�l��،bZ��Q�X:��� �q��.�R~h��J��$�������Ӹ��&�V�((���N����Ƚ7��6'���8<{Y;���m���V���s��3� K�B��_�(��<\���t��)�]����:mf�1�`��k�	@�z�ˤ�U��������3�� ]kV����j.B�t�'Y�.�g�[�!���E� m�~W} p��{�ƕ5�B��z����{�2��]�w��	���Gt4 vRb�2O�@�J�`b�q���7�C��|�
[-���.,��'�9�o�l�}�*C���N���� x	�(ˑ柗<L���O
�Q����Gc�
�ܑ��{E������AkF��Q��v�1�	F�HG�ꐻ��2��ސhy^�Bk	Qsk�	�c�������ym�gH`��|{f[L������)0G ���#GaH�Tw�"���'%�,X̓��r��g;��u��c�	q>���<�����Z�a6|�C-5ɉs诰�ch�$��k���؉'o+a��P��"��06�Y]�k�Gi����U���n�C���eN���JFVV��y�(��R�u��J[�ҿ��Hڲr�;U�A��>�=��DH��_��U23�8{�l�xE�5h����K�[���a�4��F�*ΜyJ���J'@.����C�`j�/�j���4E�C�b���t_�ͱM��gii�G�����l!7�P1
����������2�nA~�H���p��t�����z���J�f��r���t�bt���؛�����*4�e�R	I�9�g�����ϰ���Ɣ1��n?,��.��A��tC�Ё�waE�Z4+Ɋ�Oۑu������D���>_�y���8:luf%�'ޏ99##��nE>���韟�_��%c+:���Gws'.���6�֡a�1@n,CLǈ�=������2В��H�:+U����ٿ]��3u��}�"��t�[L�����H��ח��`߄�U��}���1w��`�	y�r|�,���� �g�����)�t�����n3i+�wu����)ܺ��,; k��F��_Y^���	�~˘�r��q�ss�ԋ�^�s"�cC�B��t|��|��砼���=2�f�f�01�7+��}�i�Bo�0���#�S�.�2��]��g���0i=��r��ʺ��x��l��orUP6���{��ed�����Z�Z"�lpT]*��h�%0�SERX����H�ԘG�]���X�������d��U�� 	��N�����7��`c5h=�k��uoÞ@{����r���w��6$���� ��;Zi���i"'�B�����_����@Җ���.�7/��.�teN	ک�;��~�=(gːk���\�&���F�rM���?lߨ;�|[7�JS���@.���b<Ǜ�F�����ԅV����ۿ&��h
ff��٧P'�_�	���aJ�ªiB�>��A�n�`NBB��i�r��$�J�'�ן����?��I�~@K�g���WO�p�k���h��H���������1^���5�,��H�_W�n8��|���u/1w}����%�������E�f��z�����u����=:h�q��C��WB���.s\�Q^�qڗ��4uM4'���jɤr����Lc��|���v�m�&��2Q���ˊms7
G���.��Ձ$�9��q�vf�bo�4�Lò�����h%I���3�b���*jr�u��w�����s�Q��w�0$���|�|��1�U�dpI8;F������}k �~q��w�B���J/���٦�c�Pჩ!	/H�;m�6�3�h�m]�[��$t[�nd�v�lux�k�	���~�*�\���n��3aj��\���"GV��d%�o���Oi��U���l�J[|M��#�<(��i,�
gğ��{	hS��DV�a����� ����$k�lEJ�uy�(��">�ޞ���-V�]�5`��VG��9ͮ{l
2��t�t��z�8�;[�i�a9�s��ݢ������mٮ�����Yܼ��`e�F:��&Y�_���7D	�j���n�d v�2�ek'�d��nʃ��
�B:�H�ɵ���������6� �;?[9����S�W��CJ() Z���T�Ƒ�v�Vv���%#��l���^\_%h����'d�9#�2���fk)��ј�$(~d����_��>�M��=���v��ܯ�&t���8�Z���Q��g��1�n�;_���A�;�M;�^L�xkx�=L�p���+ubj{r��l��C+�2n0S�!R�'6�.��Aqh��t�z�� YMQN�ʢ�a7�jx	��M�ẩ�^�����Q�m3ubO��Fz�GL
Դ>�J5���V�̀.0�m�3�A��}/�	��@�	<�t�S
�ց%��U .���t�4��3hxrB��''�j�,B����T{k�f�#T�;��s*��mP䐄Lr�d�xY:�z��,��m��dJ7\k�0�-��(%���pF[�]�A�w����q1I~�B���X�lȵ����*g��9q��Hұ��P�4g)g?u��M �6�H�.���H��Ѥ��IG{�+�TKw-��N���K�����1�U����Y屨��7M���y��#sNq��.[\Kl��ە�J_�2�6�讝:�N�7A�a����琼�)�(d,�[���H�A��Y�5B��@�tI�d���w�>7����<�"�}���SM5�C��P}���?���Rmtz	[���e���3�ۤ& r����Y�? �~�Ng�؀`Z���'��z�8��&�Y[o(7�R�qms!��p��S(V��u����~,*��>��'���M`H�=񫳓���4�QD��*Ve��|3�	O���R-�:!~��Ѻ�k���t�n��SR�}���=��zB��}���4��X �-P��'�/�cj�G�����D������{�����bq�q�-�2����S��<���XK�* �.���w ?��zM!�JE������(^�A�!l�Z��¦g�ǯ�? �d��:����P����͇6�ޖ���N�`Mt�Rba���+`j%�@"��}#B�(�ZG5�)��;�{mR-���VKȿ,�Q5d+&�S��\A��/�z�������5�l�-���Yo4Nrc��7n㶺��jX� �=�`����� Eq��z���w��}��/��h1ٗ�k���"?��/"�2c�vs�I��F��ڒV��I1n� ���̶ (&�v�ps��?6����)&�SS[��*���
��z�J�]����"ճ!,�_��2��uk��O�dK:.���:��PA�l�ҡ���T�\ȢB�j'����n N��u����e��;��թ6*2�$�|r�EJ�ޣ�$_���جI�t #���R1����[gB�ʹ�,4����{WC�E+�϶G!4a���8��ɳJ�`0AN�;&D_�1�J��a=�����u���t��
���)B�����~��s�tD� ^� �KnMV�����(��A1�?�M�S�_+�0�#k|��]b���fYQ8�ԉպW���Z�!�^�) ��h_�PXܨ�cт�:n[?���c��hi�.P���5͞}g��F"z}v�6��UC�P���Q�VEʩ�+Q���[&A#8��hRrÚC5��z�@~�g�7������KL��a&��
x��w���l�$�f0WX��*�	���М�P�:-�q�+�UĨ8�R����2�Z�<��ެx���kؒP�6��a=��^z"i^U��rNt�����ZRD@�� B~��µ0����8c�jm�9�!�:Jo��;�eG�2s���|�q�<�Ӎ��C��XL<kk�&�_�����`���N�ʐ��:�,�]Eɯ�Π�.��׳ɓ¦�r�d%t7�����|q����.�B���%q�h��� u�/a� �g�ֻ� ���3�n>�P�xO����dG,Ei��Eq,~��mu����	E��D^�EJk��P�Ĥ0��ч���թq�9~ߑ���5G��TGK yۃ������06���(����^یF��E�wʷ�)���(����F`�?�
�4&�k(ԉ"l�"�R�⦻�V��G��_�&ʇ/��n��YF��\�\͋;�j8F�|�����K�7�� ��}�4ժ��Cl�����)М��Sv�Y�����Q�Y5W�kĥ�U��-�0�����q��&Գc����T���ъ�A��tU!t��w/�.Y�9ڦ�]'�:��;7Qj��#��e�����c"'[8�G�! �?mg�F�^��%������S�ٳh�I����5&�Y3 ��:o/���I�m�~)�,��%�� �`��X>��%�W}�1 u#ڶ^��+��JM�� =r���-? .s��Fb'|6�����P�d�/��X��4�3}�W�
ђ]����8��J�`�����i�W�cԬ�S��Y���)����lG/i�F�����2�D�W�Ώ�惣�10�Y���`I�w���CF�j��o; ��9P�r�(�=~�Z��|��O���^ޝ�_@O��j��/��ς�P�*�x�|"o�CGf�@)�.fq�H��Zh?��s��+�����-i�M�Gcr���Ņ���	� ��)P|�4`E.й�`l�P�"�v���K�Y �x����R���ۄʛ���ͳ��q��؎��N�!��x���v������E���[Z�I�x��}h���?ܝ��R������_���E��[�����;����>���c�6)���@,#�Nϫ�t�Ȓ��j��\^�Z��u������gғs���@�� �NB��bQ��ZK�oo$�4�I7Pdʃ�ޫc��w�,M�����TL�K��fY՝�E�U6�`��?�p"]�����m�� �ìޘ-!�~����ɦ��`�.O�a��bȂ��d>"�n���=�?�Cdd���N},�)�;g"����:���l7L2k��剧���Uf�N�"�耴�V������t�l1�1Q��9��H��BmO��{�ƳўA{��:i�	���If)~$o��(�Q�Q;US��"E�ջ9����ހ�r�!+�.�JͲS�Z������[_e�'�3"�L	��K���B���Ұ�rE]u;bya�dȇ��"��������v8	cgW>G۲�IphS�Oz�\��t��ȻmC���j{ʴzu�^��2�sƜ�{פ���E������$W��n��J���^]*֘Ü��H��8��ථ� K'ol�j����:�}n�{ FZ�g
�F,�!��j��s=rS���ۯ��s��)�W=^��<�9i�~�xq�: ���&�I�0,���E9_z�iFl98}��![[��)�����'��qt����I��ܢz��o�osL��\�yeW�R8e�z0˶U�t��7���l���1���t��U_���.Alf�0�t
#�\�Bf�P���I�`��d-��e�k�l�^�a��rt{#�������?cK�e�~�W�l-���А��cW������ے��Ƣ�PG�U�̚��_a���X���qK�؉0O��1�{�Ե�2�3w����++sEu�a�FB�)�uX?M9�q>w���
���&J~�x7��eXG���ȸ��Y$���]��^��М�nƠa�!���b�4��	�B�偮�N}�ږ����ӾkLQ��b.����A��գ��,�O��r��`�>zh�m/�0�xr$��J H3y�����4���Åҷ"+3m�7!V���PKf6n	˨�]2baOs_oo� �������<��ڨ	ƞ��Jn�t��,�o�L��k!e�����l(�WZj~/�cDk���8P�F@��&�c�Ys�����Z3M�w�wÄ�?n���'V��s`��Qs63a^�k��(�"Nj֋(����ސߵ7Tk/ڿ~ː.Un���F0���S��,��z*̉���~&G�ѯBb%�V���$%�KwN;��S��&Ĕ�����.PT�V�;�vmf�Y19�,it>41����e�Lq�]fN�C��1�O"��*3��R�E���.�刾�UΥq���]�ZC>�����`h@Y�Лq'�:,Pm����Ŵ�/˕h�
�k#�=� �[��!������54�����T�����Ԁ���>��U$�R̵k��410�w3�p��p�Nv��ӍwO�ߟ���֢�hYT>�q�����̴;��H�E���ͥ<xc��KKn<>��<�VG�đ>@ Z�=e�y���~��a�l&y�8	�����Γ�hui�7�QeH��!��H��@1�Hv�s�B��7�|���	"�\vHx�3��y���l�jJ+��[m�k�XD��{�j�.x�ԍJ�vB*K�GU�l_ ��c�������/��� �u�l���a`�]�����w��`r�X<_����$/�i�9�ٲ�s°��C��b�9�ҧg8[��6�.���$�UX�$��,�i����C5������
 v�-J��
�K���������1��!Z��|�/�|c�2~�[�M`\mS�8r��{x�Vi�:-� v!��J�`���C�ih�]ܿ�1\��F��X\��@TP}��3�M�f�}D�l;����	j��PS�]=���]Q�J��QԆ��~��:1+p��E��O������ުc��xY�R�XI���;��#�
�ľ�U��;�@8C{<��4�*%�1�(ֱz!���O*���'Q<�+&EX����G�2�@�`m�c��d�DG�K1���.�	cc���GR�Hvn�_����x<�Ӯ-n���/������P��X1�/�����|�%2��V�k�-��?qX9���>�߈�.L[���j.��x&9�����p�{v#=h��u֒f��|�*��j���Lb[N0�9ؽxө��,z ;��x5�F�f�^Ա��X,�9��/ܾ�'� }~ر��Bd},�2��o���s�1���	<OD���L��*��^?���>]�	���C�X���%�R�}�����}��I���E����H���Y���U�:}Vb�9�a,Y\. f/��zؿ�ת�K�����B��r��Zp �~wt&�1�-��81�:��m{�x˾0�#@Ḡ}^�S�J������� n3�z���;�w)��c
������nr,8�Rh @���4�(R~��Fl7��vu��Id�t`4�����m�ߝ�w%�[��a<�:���u,U	�`)ΈChF���J��+����?$�7���򃹡����p=��tt?����JQ+ǽ��q��ڄ��������ٺN��~6AB�~.�4SPI�W{k- ���+˹���*�����L+��S�������:��>Y��gB��0�]i�k
c7ؚ3;��\�|Ѐ�!׹��%}Ip7��#�ɪ�9g;ag >/�U_B&�c����!Sy��9�<;�־@`����[�LS��b�U��a%5V5$��+`�g����7��w�ͶI�jC4����Hא$~G�7�V�k��1v�B��*�=�D��[�q���_���19����3��;�7A�Lܳ�-�ị�}$N���F��0���I(�'E��r+����:�߼��1�_�%����I:Kq��Pv��k}�oz�5�~�k�2�-�J�_��{-5���ү3�BN	��Ağ�Q\p��������h��X��2gU�d���[y��3��}V��AL9i�&����%��v�~丼�ف�a�Q� U��� �����X�9ZS����5�w����7��EQ�ɔ�������TO�?��]���*\j��	�lEaY��B�8HI�u�fvd4�%��)������#�l�=���X
����l��0���gr/z�I�.6�/�q{2dߡ�.%�G��v]Ƥ�q3ڇ��x׊�x�ڿ]S|yMڊub(�'"�\��(@g#	���[kq�j�d��LY�'�1!u�������C�T����ا,��$�tyg�ad�]�}�������3��BU��?��V��J}�a��Z�$�f��eOÎD��S8�E�D���Xj	�peG49��)�]�z"*q�O5U�c�����F�����O?8ȼcҩ���ϸ���x"����[awc�̏����e���y]2�p�v�W�.���¾e��WD�V�b��ڦ47�B�2Q}y�$�v�a�k#ٲ
�������D4)�4����6�M�v��h���QQs}+�;3-�#��7{���I�B����]*��-����$��h�u(�����/O�0�Y3(��R!kn���0��r�j��)��ޠ�~T�@����
}l����`��_�ڿ��Hy�p�|�o)����` A��U���f���)�]\ ,G��S׍��X��ڀ�Y�Ic��g��U]�f�5=��1P���#A�cF����j4������u��UgE��[!Th@�;�Ԝz����%��5K� �4�?=N�s���E�e��o�N�uUω-PA�ёxo�b���)�;Ϡ��kx���m�@�)�o�䁑u�m�
~��!q�x�]��Eͧh}�;�s(�K���TUș�L5y��R�rl��S6%BO����\�v�$�	�sSO�6�j�^�q�
2H�$����\yhS��3�U��Ȫ�4�U����4�3�F;Y,˻%$������΅�#ש��!r��i8���� �yTj�W%J����`<}�P��T���3N�k��I��I� /püZ�[2ׅ�c6���o�m�ׇ\�$�UD���A�T�����'���}���Z۔������f�Vjp�����d�d\�c��_ؙ���3�A���Sؑ���g�z��tR�e��:�K����-�U� ո�΍o
?1R��紗7�B��nS�-s��t�͵�i� ��}�dE��:�%����#L�5&�����7����n����-�֤ޛ{8�U#0�jDV�ƘШ���Z�rg.���-���:&;�Em7a��_ �ɼ�R(Ӂ4�u�6)s�&�냝�GR��� "��"�D���ۨjfgH���ژH�A����9-*��a�`���k�j�]�އ��[+�C���Gk6J�Zd8���Be-��y�5�('�G1/�p'b�1xd��kV��B��ҷ'��_Ŋ�8͆MaT9[
6�\D،w߄��/IdT~�̹�3��a�������x�������y�$_Ob��T�;)gXJ��	5;�["Sg�'` P�k�v�碢W_��A��ղ�%Z���饁���42@aB�]Ϗ�Oh�k㘯��N)n�n�B�IHG�*M#Q�}�r(ٚ�4���:��v��K�  o,˃vs����գ���v��da��6O)��+�o��B�|�R u�I�,3r�����Ҟ�=}�5J}�w~I�Ӑ��}��3�3��k7R�J1
���,�Yv{�K\V�ҥ��8R�ך���m	��2�O'َa�h��/��׆�!�U/�t���{{L��}!�6*���"F���܃e��뫹X��7q�8�S��D������MRS����p�=}��`Jo�n���zc�?���h��x8X]�K$-Y Ջ(�T91���Ar�i�9u6/RPI����wұ�� �Rv]W��X���2P[7�m�����^:\m>�^���0�)���Ie?���07_ȗi1IB��r�K�K��č۳��<`�R��_H�D�� �>>;iې̈ ��(*Mo�Y�UJn����Vt�8w�H>g������6�J�`� ��|q	�\��"C���7�Ԉ�c���WP�j�ֶ̚�A�V)���T}�c_�� mM)��H:�e\Ҕ�u+�-����J����(d�&k��)�}�(��|s
3|}�{%�8$C���B��=B�"��:�ی��!HCP�i�UP	��S�Z�@׾C�,LF8����OY�h���>7] ���#�܇X��P4���u�i�B��P�E+uq�i5��ތ%
��������A���i���D:_�[7�h�o�z0���G�����#M�`.��%�p��R��$`�텫R�#�ޟ!���ں��,�w1v�{6�Ɇ�� [��$�{�=���1�:���7y�S�i}�-����[h֏���f���3��5���߁Y��7^��*��M��	3m�i��IGZ������-��|<�Ŗ�o��i�෹�oԜxXf�A=��G�5,�Ň����"<�L���aԏ�����Ҕ\p#�5p5�=���] ̓#J��qS��.
j�T�U�Z���ɾt��E4at���%��iA�^A|��b?%�0��=b�j�����\��3>�?Z�R�3�<$����5sr�Y�%���˹tDJ��[
�wB\��ұSw~�+B�����{M:D�&u�Ӄ^�X���d���3R�M��B�s����NѴ�ڱ�!�*�I�{�#�s�g�Y��/��{��p��G�jg"{��ĤMű�W�jjD;TY���3VO2(��R��/~��$g���)}.ק���:ӸW�)�X׳�}����:�:�kYi`[Ԫ�`���t��-@��F �����b�M_ؿ'*�lY�J2ȼ�����ef,��9�b��^q��雖�2�����0���t)���X0!�e���+���{�+�EsG���u�S����.�(�PmEC�Z�>-J����HMwmAZa��:s]i]G�Ua�� ��E��b��׳�xh�s&	q��EM4������$�KL�K�o���z�����p�G��PS)��N`hN��TQ�Y��$����V�Qyx��+�_"g� �����g��;8�aW ��A�=��h�pY�����j)��&ݥT�0C�_�ࡹ\���\Uq��]��]A�a�g�<��Y�l�@��l.�=�#� Ӫ�c<}� �v��Y%r6���L�����|ޠ�����.�'�<M˛_��i�"Y���n8�źW5c��}SpJE�45�z��.A^s-���#� 7��4���m1?�haQ��������f��}n&Q�W�5�8�k- g�rW�_�Ҳ�Y��u\O�������F��a��n3�8��WP��B�y������� �*��:O����Sp��{j�8�D�V����6q8Gí֦Vܞ�o���%l`�8G@H�I�A�4s�\�
� .��N`��`�=���g�'���v���az�]���a�b��*�T0�y\]��Sή��q,��:ɊBT<��N7O�5&[�S�R�@���(�{t�	��k�P;�r�꾸$�E�`���U��e��Ǐ��4�?vӕ����}�]\WJK��3�r�M�Rj�����x��t�_ʛ��/����w�~�`��I�t�ں���h?�e4&�}�|Ȧ���ǘ�����?�헁?l�ϝ�M](ߩ'y��f\�c����zdYlV(�'�%�i�0h�y���J0w�Ke�V�δt��ߥ.��%I
��� ҷų��A��ғ�����8�	N'ʇ,}Q�N��R�&cf��B��gR�ͺ�2
X��^d�V�q/����-���J=�1�57��t���[�.��J7����*�r���2:��Kve=�(C�>1���@��Y�q�t�av_H��5`�*�ծ\��պ�E��w�$�f�a����/2���x���gK=c�|Tq6dHn�D)�ca��{��WJ�Q���r$)�(N��f�0�Y>L��|��t�������m0��m��1���(:�9���������h��|�$!�P�g�'K�f��"g8
;24k���`�@�)"e�rI�@�.��U����5A��t� $bjÖڦP.�����O;���H6a�. zJ�l���~�����k�sˢ�JNh���PI���c{�Ig�!m�F���"�.L��c�=��D��_C���m�8�����/�&�����3E�q�h^�]��'�wy�eX,�t����� u�_0%�,~26͗59j�i-S�#�pϧ�+���]yY"�t�}�O��ć8G�5 ������ڣ�5���]��<��9�垫�չ4��10��Ԝ���k�!�р�)��?7���۟�)���m��i��4������p�:{ܾ�T���+}�3�	v���moɚ�tN?c�=a�,Ѐ��9�;�X�i��3S��"��~��rҏ���
�+O�"?jMN���cr���p���[L��j	���_�tx��P��k�y¡�9Lm%��2e�t�ez��E�/�gX��u�ɟĨIkM�(q�/-:�НY�Q�o�ʵR���7�/��w+"j�����`���䓦-DWS_j3��ä`�ӻ��s�w�v�g�����NIh�%�|�&՚[:j��R��v�{`1��֙�DJ<7�B>*x`�/��z�A/^,�`o����&��|Ubr�c%�#���(x��<%�9�\8)�����Ԃ���5gR[��#�����9���W�]��� ?_o�J61"�ߴ	(�̂�Uh'z<�������5zIX٬���TAbM\$U�E��e��(ޒa\������;����+����p��y��aM�2�#��C��;[��(� ��g�ne�ELH�r:}q"<�{��E�Þ�T!ϼ0�@|o�""�;���J���4ż,���U ��
�8���DSG�̱D���c�Y#�������������𝑒�2ǥ��c��
�;1H�=T�p����v�%�mӯp׆��Kp�+ʮ�?���n�����A����ó�O��W�\��'�!,ƥ��<r�K�ceu;���	.������=�.m3d��0U���Frc�9�io�u�r,L��ѯ��^�`cl�(�{/< X`aDK!_����s?��P�����}���͂�K��V�侧����6��D���@Q2Hv#�`q!*�-4�����n�����ޛ9�L�}�(~���RL�s;�{�R}%���2��C�
{�Jh/
1�?�0GiA��#�Ě��Ud0���ϓ��,W����şʙˣ!ٲa��#H"E}�\9>J��u߸ópR��� +µ��Z�M��<�:�f���A�цs�����th���i��!��r���G-��=��d����[�b���{I5[�(;���Sx������c�TwF�$�F��[2�3�`b����	w�PwiIDi�<���{l�^@<A����k�q�9x�&��G�E��D&5�w��&�Ĳ�-t��˯�rX�����p�/l�ep�fR�9�S�pP�O��V5�_�#��ä.�����E����؀��!�8k��};�]���e��u�am�z��ŋ�P���s�*LgG�����5xmFk�Ŕ��/�8u�7�B�g��f���=�ݰ]����%ˇ	�Бi Sw�R�SMٟ���x��]���P���N&�9h���m����=�#ش�7�8m��E�bO*���#���4	TJ�TQQ�T:����+)��<v~�V7[<�z1���}�9�y������!HO��6~ߵ��o�	��d�/�8�� �V��9��0Da�1��/m��a�S��LnP�G���bi91һ��vf��｜�h����*c(~В�M���J}UW��3���8��p�9J2�ݺ�W�U^���ʧ\���X��K��e��������g��שJ�����ي��J�g��^Z�Ac�uy˸e,k���ޑ�6ň�JJ
9�2��x�0?�rI�iw�=���;�M��tUG3��V��Fk����f$��m����8y�	�����9�g�`Y�ŉ���ʠ��ɵ�����U�(�ڦAB]\P� ���Aɺ�W���~a��w@����"�b���6���t=E*J�����DWq��;�a?�ov�˒8����}��Ҁ�b��핈��
+�l~u�tN�=��趧�3;���3��=q�����¢<���K֥RLm��&3������J����꤉m2ruSu�,��D}Rm,� J��`��6E%���.�g?��(�����2��L�ex��
�6�W�&�
�݌�6�T��5`�`D�k$!Ғk�G��+��B��j�Eq��e%r�g�4YWyZ�:����]���^g�4|_K�ę6�k���H3mͲ3>L i�G��<�{�p�����	��G���>]\�Zڛ��:�l�[����/��ӂp������T�ؚJzA'>~@3�yay��L!DFٻ& �q�k]LV�aã��ۦ%��V8����<�,�%a�UtqN^m�]J }�&SS5�|4�����-?�P�((��8d߳�PQ�'����&a�,�]Z���(r�B)e/I>9�RWy�vù���m�"��E�N�Ό�+�p  '�Ә]]s�f�H����`�H�Au_��*��=��	Lm��*q��O��4J�smV�9��%ngg��Q=� �ɺ�9���TS/�OVȝG�]����CH_l4f�Iu�@8��+{"���:���օ�����o�myJhy��X�cu����Iz��Z���B���x
rw����01(~_#iU.F��ן-#2Mk&]	#�������j���@��w8����mo�Y�����l���3�mz�� ���|S�� ���PD��F�T]�����0�~(�mf�Z��[6��^Y��u"���T�գrLGʹ���t/r=>f'k���^V߃Ѵ���_��]3���:	q�^o?B�&
@���֋�HI�����n�g����֌Iw�-Y�i�u3�̅y��������8'����Ҧ,�_���K
>��"D0��@�*AM�U������zƃ���SrF؛��s�鳱H�f�,ޥǅ-����߃��2���_��~̳���}����ƌ��)�O���̩Iө�ݮ���,��3,u�	M/�\���-R w��c�*�`�hv�c��������&j�>�*���}[�C�#���!�*C��I�J6�\9�'ܻ���M3�������}`	�j�u/��,R� R��e�
+�&�My4|�L��32��gc�/�|�Z���lƾӍ�n�8�9�	��l*��ܑ#0�A��=�_v�_���i�K�Lz�����L[��L�	��9go��C~�p�$H{]WLʫM��c6i���C��׷j�ՙ�D_tN4�{�Z�����'<#�g"*�`
5W���V�0J�}�I&���"�3&C�<�b�l��N�׀7�2�}�d�k�m�+�ܧ߰�z�|L�+R�]�nXW1�o%dIx��/��Q�KǛ���ʴn�g�J�V�%{e����Zz�hhg9;�`,<�.[�#r�M�'�x�����@Ұ��R���3��QH-J��E�gK�}q♅J��Sh,֥���<�<��[S�b��i�{���_�uT�J
0�����-����l��Hiʄ.��o�����)$�P�c���rvlש��X@��AA���I���1���ɲ��?GꝪ�e蹟�x�>���;$��.�-� X:�32��,��2N+�w�qP��L�a�AT�M-������TC3��|C�}�Dl��:�"�{iQ�0�:K!�to�$'��}���FF5��,6����L���-wn�x�S�E&4��z�����|L��'I���F��	@��w���(�����C(�eOY�N�q#�&=������y$��2�M�IIל�s��#"�N��	��-�y6]foC�V�Q{Jz xP,Wb9r+nr�wQ�Z�2�H-��c����9�������Ci8�!z5~���PT��ʊ��4�1D�'�k�4�N�ʅ��u��2�3�F�tI�h|*x?\
6cn��p���[�8��l90^�t'��~Z�Em�-4�=�g�8�[�4<�����4�A��uxYQ�m�7�Pq�]��ϰ���<蛘\�x�y���cb��R�5_LH�]�F��m&�
k��Ы��7�����]�sO��1zo��H��yy�B n�j��kb�������1����˙��V�C`�j_���� ���VY�!��������eq6�>#y��2=��J�:~�>�p׽a�� ����΀.=UC���) +�I"�9�:V�CnKƔ�L/#k�<�v$R���4��4(���iL1o�hD���^nn����u�52����k�<���P�l#Gm⵻�ro����^z�Yz92qj F�!6�k��3��+�UQ�H��gג�,`b.x��z��lb�>��X�p.�i EJ>(�`O�~��:`�٣n�Xn�h��,J>tsqOSqԾ��c��;��� 9�C\�	��n3��'Z�2oГ�ڨ�~�oy�rsY#H,�{����F�!�N��}�Q�ʝ���e��S�k!�^�_ze���tV�"}�G�"C(��NG����w���D�����^8����S�#t�+��#A�`�'��UQ�I���l���_�h>��t������*�����(3tGY92��T��Jmh�Mp����'�J��o"*mQ>�N���d70^�8��R|!��w�='ܦ�8c4�������$�A���P�*�A/�:���i;��Do�y~prM�N/��%+g�/�+[� F�YnYT'?Y�f�~#����8�r�ڪ�3	������F���U�HZK>||����{onf����{���e����n��]܃]� � g=��*4�ka�UsT�tpc�˭�!ny��	�¶v}�Hq�N��/���ʱ(�z�S<��W����m�����:G��y����u�\g�FN�nZI	�QV�E�.���>��vT|��+y4)�ָn����,�K՘1�&N�K���I��s���鞍(k�"H���v���h=�L(������E�!�NHݟ6PnG�g�޾�����&O;���9}Ϭ��`<2g%��Z�7<_1Σ���a[��8QTp�u
�[�i� �<��	��W��w�c��p�{��6ipʲ�'�~���̔��@C���a�;e� w��G���(`��o�9S��"R�Q~+G$�q��p����fg�I�1ѺH�,7���AX�0<x����?�20"��8��]�ұ�����e�	4ߙ�GޤR��m>	��64
�5���eN
򮜳D;n�E�lͩ�-����!���@��^PJ�%A:���p�y�Æ���e��9Q�2�y@'K�����{پ����.?�d����}���1���H�%���-V�Mo��S��V_(�>��ݤ����x˒�ܰ����x�Y�*�����d�/Qa��ll��ᔈ�lx���&�ǒ�ɄC)����[٣��6�.!�y-�,u8�fǎsg�f�����}���A�A
��%�p1�Z$�����-��h�g�����7��>�H�( ���m�>�-�3&��U�uR��Ps�ͷ�kC wh��vQ;{j�������̷��OX#S���-��e	q��٤�Z��2 s�������F8��:o����N��1k��UZ$��j�5I��J	"�$c/�n�DP9�j�R���ӊ%�G���ޜC,�7������(�jf㓓�*��¦Ӂ$���wL�;!J�^f�U%KfKzz�,���s{Sf���&�B����A�e���]�Ë,L0���ݫ-��S�?q,��jy�۾�q��Fu0�5����ـ��G��7����bf�*$�:�W�������6�o�[��o�%�!�@G��]4��K��b�J%5���6�_�bJM�e�����Q| �����R�N�bZ���e4�h���)�2��+T�:��0�(y�x��xZl�z��*���SB�Z��Z'��O|�9�����%�0Kmϴ/�9���� +���~�������*a趶��~�(b;<�(f	�!8w�J�J�9���7],%�.��ӣ�̗�k��c�kt�`�&�9� �&���LÚ��¼r�c��-�t�:�/R�d('�t�����-�4�
������F�!�����V��&�ܴnTwR�����ҡ�u�3�i��P�uj��_��,��9��o��5ᨕ�������*���j�O��#�����#��S q��c�.ɴ�ip-ܛ��e�f�+��J�@�ӵ�׾�_�Ē>�NV�q��Ғc�1(��yK��J� ,v��Ъ���}���҆R�JJ�s�.}bP���x����e���4={��JyT �����׫p���o�
��������ZbB��	HHx����Te��>�"r��d�Y��0�]F@~��������R6�S���L�|��j��Mr�1����9a�]gW��%� �dP,�>�\p�gS��4ۍs��S�B：��F��;��&���lv�L_����x��6�7�1�_fkz�MXk�j�G<3M�]���V����$���Iw/�8�rzv�������f�H��As�^�$(��l	�u�X��}�sR��<�JE7v��llV�g�[=���1�$�+F���Ha�8����J���.�yU�e�&� ��τȴ$[�s���4��ȑK��5Q����kB��2,�:;G�� ʂ\�a��ﭒ��:�߯�c-y�:]�r�C�B���b�.�{�e=@#������ѩD9�K %��B�b#
ܾV�~S�K�N��0AT����N١��{�e�9g?\��qG/41�'2wAk���Ů�7M���n������b��hҍ/�1�쏾�D��8n��9G����գ{�6�W��e�%��+�Z�E��&Ad�F#��⍗����Hk#�ד����&�Il�E��s��b�V���G�i��~>)͸��>��o���O�,�\��H�84FV_�3z�J���Hꡁ��'� ㆕J8��B`nr�U���О����a��0x?���r�]����AuddH�<����cd��h��!����6�2W{�}����؟ٟ��;A���;(�����]Ёk"@��1�i� t퐠��a���&7�+�3����0R)�?�T��� 0���\�'��r���А����>�����
ԭw��/��5�~7���I �J�1J���`����d$ۀ�f0Y���sc|���f��m�dE��=��Z�OG*�˺�V�{EG�`�dJ^��?����$��Ł�%��0[��|<��eG���8���!�A��L�&�cx͇	��j����R�����@��k��j��u+M��v>/����4�/�	#�N�D55�Ʒ�S�4�s��V�(ZX؀�Oe_�f��;u\�ֻn'v}4N��$���j�l}�a�x@ֶ�
a�)�0��tg��T ��&��Q;�&���sKB�Hs��W8娆���ڗ��dG�q��+�+�o�B�3b���خ�^��\@���J>�W�.#qJ�ߦ��$�u5�m6���Av9Ţ�6� T���T�߂����x�!.�)4
�62>L��r��hwP�,ݪ�
}%��cG_�5���l�۫I��bB������=�]��O�͈X}�Xs|��㺺S��.�Y�Q���	�ȤJڵ1���>��Q�fOX� \4��"�Ϡ�9��t�l��5��\y�[~[J�1[f�0?�N���e5��N?ol����}A�����H���yB~2���V�q�k�,[�Dk�ό���s��O�����ӕ	^ѹ��U�1_�}f�{�{�G�¶aq&e��ߵ:@䆓/L&��羊0v�T>J�����_�&��RTtm�l�	���b������g�rdI]��< �~=�z�"u�4b�"�[r��@-��ɠ�I�A�*���mcV�2���h�qV���	H�N��V�8�)����Ii~��
����Ư�8��B�a����~��0Xˀ�-���vB�6k��1u�ӇΠU��0;�v��%�ؔ1*�D���yq�wJx?Ѭ�Pt7x�����F){��1��y�U�m�[0���Z����0B����q��i
����6��J-�a& .S�"$b��@���M�X��%e�l٠�n����&�2����4�'�[��~|���
ن����P ���]�) 1�Q��F��m)�������H
�	C$Ͻ����OG��f�#,:o�Q�Y��`���&����G��6re&����u����Sbn]�����{���U�z��`��oS�H���C!��sEN0．k�/��=��]AQ^z�ɂ�ޝߕ2��l���piD��)�����Y����d@�7��VG�rQ>I�C
'1.��[$-���"�b�ZR@���9U(#��)	>�k��#&u���3�S����oDQ����u��<�_��躖]�Y���m����|ާY��'��+85������P^п�L�aYac�5�2�p�6�=(2�d��\���v.v����Vp--��+�u϶��e��=hzZ���K^����k��y�����{��d1}�3y&Qu����<GE	�C77�M�P�Ɛ2�5S�2�>���'WS�s6�=��W�B@d�{W�];3\:�?�E{�?M;:�
��ڥtCOX�Zz�$���7p��$";lԄ�7^�>?�z6hui6�,�~�f�C0�O���������٥ S�]:����������r�/�C���Or�U���\�}W�m!�TWp�8���,d�ҝ�G���E����9�(�����Z:
�~���&+�g�x�v��zKS�P˔�S�3#A�f��j�"~d��G��6!cag����.�{�D�.��ò-�4�+y�֫�Ld!�ڭ�5mN:��v�g�ݕL*�r��uUU9xu�]+�xl�1d��F&]���b�Ԥ<�GGA������k�*���;9�T�x��z�qy�Il�&媰����`	��̍N��#@^}����b�)xBᎌ#��Ł�KN�sQ��93/�MY��s����3q"�g��3�
�'Y�uvb���B��yJ�!��#DJ��뙱����Ď8K�J����zNE��ڭ�־�@�˞���,ny��aVo��<ľ��オ�oܽ��fk�����.����/�M���(�L�j�1-ӹ;���+��1O�>$��Z�o8�v�e1<����
P^>�o0�MIʏ}T��!��G�hD��۠��`�
hӱ
��+��/�1�PWR�cd�R�\�EL8�J�du�>�y�\~�i�aN#��'=��������u5���X�����Ȝ�_냋���4��<e��O�����L?@7 �sL�#��b���}�O���ڰ��ug�R�2R t�4�#
{#��<�AM(�yV0b\��3�W�;��o���N�Z��!�An����|��6�7�c����)W�Xɬ�0�d�Gi��s������ ݶ�s6�di��X�1�������+kl�A�4���f�`laV_l��X?�c�q�6�P�K���r��8)#��W�#4K�.N�N6��q�M�<ǋn3���9E��{�#ϖ	��-��K�V�W�Y�X(Ft�x�=$�%	}fMfmJs�=��P+��6�Nh���]>j�Fꈆ��q%)3��5�Â���]C�)d��/�����v���l�������%t�m��.�t��l��f�r�p{�o;��"�3U<Ds%��sί+6��3�[e�{F%�'�b�u��}� ���~{��Y������<2�7�v�I��v�a&ey$p�>-~O��;)N��i�N_��	�C�_��H!_ѱ����p�f8e[��{�����*�[w2�c�cj���EZ�b���m�E������-xU��;d����9�f�*B�s��e��`��$��
r��d�P󯛬'G�1�V��p!���e=w���[>���p�&F�ŦЕ��:�/��g�/�Ew�_�jU�$�3�""�Ԏw=�=��;��{}���qL����Β�O�5\�D��M��0~��a�8΢`�V���N��׏�o��j��A�wN��U��N#B(P:����GQ�X���g�,0���>�S?	�h@|OG��0�E�Oе�ݲ��N�	��<��V-�5 �zv ��j0Ε�k�P���s��e�&^�D�X���nj��9İNF���:�|�Ј��T�[�;�l��9�4w�Y���t�#x��?����咫Ck�S���9��v����Q��}"�lx�1���%���z�%�o���Gv��؆����8�!Vf��\,���eu��<�����V��Z�MV﫦���w��Օ~���Д�M����� K�;)O��*��S!5��H�K�d���/�'b�]��h:kI��@�����ݚvJwQ�&6y�x��7a	k����5к��r}�Cu�T�Q�y�'6v*DY�0�B�8��c�@F;@���3���0�<P9��-6�QY$�ų{���猍�Q�N���JF�c ��8ɣc�^%� |�������˅� ��z_�Mj��ݛ"C�6jx7�=��88����o�̆(��G��$ߙ�t�R�!�J�9�I�u!�a���J��Е&����yw�S��*����]��Lk��r�� ���d�����F�n|����7ڮU���7��k����G�r����\���_`�b�����-C����e���~�m���)�|UU�K6��a ��5�[0^[sjϳg{�����\��o��P=�z�{Km��6���6��2W�ݹ�`�/��z8~�> ��ۖ-.�l��ڼql��^�����Dm:#D� b$+����sJ��5/ݩ���?(�鲿�������'1�B7p�C3v�ЫȪ�h��aw���h�r)�5�ۮv�T����>
��O���^���WF�*�&�o���O��R���`�W��[:$0��		��L,ȳ���\�m�Ͽ�H#1��*Ʀ��(>�S��7{�b����4���hJEG�(�-b�Si���;�f;�j ,���@��uD�R�s��*�;$P!�`�%�3�q�3�g)Iz�[/TH6!Fr��Ls]8����
�`��g�r���a�u�1Hj@ᬩ����<xJ0��lj����k!�^)���SR�S `,��������׿%��;s�����KB�!=��)'�/��O�}�k9���E3��& �
P���f1�F�WV��ޢ��$�J��Mvt��#�FXZ?��1%)��3t���R�j����� � >;	��u�F�<0����3^���M�r�>p��fȠY~E诧�	��1x�^j���.H`+�n�@�6��@�BVG�r*۔���/Y&������&�~�!e�g���]��N�d9Ͱx��N�Qji��]Υ�M �����خ�g5_�RR)��r���P�\��;��+(�� �F��Դ߇<d�l�g�;�'�)�����Tϻ)|��VN�&E��Q��Z��ɴ�x���((ү(����o:QB���Èh>9~2n0YҔtN,�*�e�	ɪX�������+l�]�����Ľ�<�ϞIe������6|�]�=�[1���눵�8Q>k����vN�[zD0��3H'~��F�����m��k��ou�������t�s�&n��%�m0{��.�2 ��ls=Y��q�{�QJf;��;K̊�����b��Ts��k.vڱf��j
x��>Y���*Vy=���⾪�9:����ƣ5;�2�=���u��UY���}���������C�߉6��W; ���]��/��]~�+�]��A89��rD(��tu�@��\Bw����	�ZK�/^�e�Ĝ�%L�㧾{�q�Uߨ �X� �ҽY��^�噴g��jLpN��_(\�@^�ti&�^�cl�8��߳h��T�=���dU<#��9��Y�8�/b ���a߈���'��59p��q/qQh�F��C�j+3�/i��c�(��Bx,Lm��E�/����F~�+f'�O�������S2OnT��:yc��\�LcY
�񟿵qJ�<.[DS�뾟KoZ����n��g�"A�vv����&�l����=s��.��k7����4�uE*�=�wɰ>F�q��
�B#�r��N8/�H6�IP�����M����ɗ����i�P8�r�]������� mU��d���gL�ॲp��e��A�L?>�w�+��4�N�s�y��K ����@>$�1U��f{0�tىn�z:���{����.��ç��W0l_��Kb�@<�&w�>��EC�,��>U��I[M��D��ύ�%�6���`�`���<�&&���~��"{�Z��Ȫri��e�Yr� �:���B}�$��j�dQ�����m��x�Rf�(Q�ɔ�>~B|�+]���WK�,P�@�E�nT|C3�m�*F�I.�l�b��$�AAP���`Ñ-����"���e�?�m�1�M���b �)�w|2N�I�Y� *� ^0�3�
h�'k��`����>������[��(�}�-���l�7l��$�NЇ_6a�wP���潟Kj��q��"��*�V�'��j�uF�S�R������:6'�@�B�d=H=+OlT�d��b~�z*D�7�<b6�.h7*H�������Z�YBĲ�4#�E6���D�]�Zס��7/���W�S��4���f��m'���&�ʓ��R��1c��ۜ�ʞR��L���p��ܶ�k}���g� 	*�uf/:��V`C��� �\��ɗ�?�DV8@X��L����Ū��>��Mh��>x\�{�e���O�婜���m �d,X�Ymr�����$�L�g�g<a�'/c'Xx ����sL��G4���w�X94')L%h�*�:7y{�d��F9�t�� ؕ��s���:�m��K� �n�#����Z����$����}5[H�#eA�!�1� -�Kѻ�_V|���&��i��Q�xt����Q柲�J/��AJ}2���:�+�6�
���Z�눌"*�s���r�����1��7�
{��Ϋ�[�9�/(,���H�G,3�/�N蚇�Ԥ +Ϭ��k�cR\�YXJE9I)���]'�3
�0�� g�>d4���W_f�}���^'�S�<(g�t;�A���n����M��x��F�l_�iwF��'�w�$@��������Z���N��i�}�X���~����K�@'��)��mCZvT��=��������(o-���k�m�Hs�΁��Wt��'���Û1����}�Vb��Qޮ�sTX�S:�V�-�3w��xp:����i;(:ג~�U��!w���0�&#3���"�|?L�u��W��U�^W7C*TЇ���hs�uS�`�	��/�~��R����׺���*�F\�HYP�Ӈ���q.e��No3�L�A�;����#�6S�(GW�9E�IL�2��J����6�G��ǂjwT�e糕
�l�W�CpK�帓�yC�]@��^R��(�}��_�vG��f���^�pp�Vn��� r�7��jj�
Z�d�����CTYA��r�͘�K�,$z9��S���c���� hJ���pT���N-�1B��c.�n޷����O ,&}�0��W׶�&������vE$�k`���ƛXQ[j�2qS����{� �~�<����!���_�9�o���P_?���ƌs;�t�r�Ts�L��:z1�B��Q��j�` �����_/��6���YcyL>�A`��=�D����>�)�`2c
A팛&�[@�{G.�HP��s9Γr�w֢-��Q&?9?%ܖ� N:�)�>JHڡKF��{���XxQ���:��N��ħ�}���R�-( �#`���9�S+R襔�n�X�ё۸�3�cwc)�:+ַ�n���F��}"#RϞ���n��+g>Z�49�ꓼF�I:
�V*I�d$�u�%3�|� �&�Z�Ӑ�O�M��Ƣ<C�OH������M��������g�?��l�#����	#�)�j`@�w�J9�xN1���r�JG�1��eY����r���ׇ�N�%f�zBb烓S�,�;�Q��#{���~���� �1�gh�3�e#���hٞ�W~�p�}��L�u�\���L��
��t����$I(�xs�N�h��6�Ӯ�ob��x�1��4�E���/һ��(�nA�qk��+�-�q�& On�g�:�ߔO���_?7�G�Õ%(�+�]���a祍�L\��q��y�Q���sӾ()����.�Yk�&��~�4f����c^�W�Q-�з��gU��E��Ί��&�8��F��.�ߟ�`����-Ɩ��n��xO���]4{����>Q���%e��g���H���ry���n}D����cj��3�����#����e�Y[������29G�`�">צ�nԌ�Yq���#T\�jN���Ў�`�FC�ƿ�*?Ą�n�ܪM�j�|L��;����QP:�;9�v�0Ki�>
���L��aխx�M���*G�R"a�ܽ,B־5�F:AA�7�M�`zXE|[j����KW�J�T�W�#8=w���	����Y�
 �K�5�}�Af���Ƕ�|V�i��^��s��eu���c\���u>�zI���w)�{�l�lZ��E�P[˗Em�	��}�S��bX��s��67���m�㙏�)-1��@.D�p̷������x��E�s��k�= A�*AI��E�*�)�M��!�2��}�
z�2*��p����u�����О�
zk_$�ㄇ�8QRkFk��j�[�1�I�` "��f�\ii�`�t]��-D:E#�O~�s����<�WǗ&#�C�]��-�PX�>2p%�Z��6�t�*�wG��\��%2��}W�\YijPZ݄�n�Y�է׵��d/�|�06��(��>��GEsJ��>���#'�rb�Ɛ&�a⥝��m�B��)MyU��h�7Z��yi#�*�%�|��C��T�#�8g��y�j�`z}^bHq�|�#P2�r���-�_+�m�c,m4��ΓLy{\]�����W]�E8��"-�	���Z�N?�Q\t�̔�O�K�h���C�0��:���#G��C�F]�)���Sj*���F'�YV�c���;��!v�ߚ����$|jzA���4��k)>�1fvy��^��nc~���MU6g��m�V�� Sbo�i�I�TщqW*VM$��ft7���y��������.�z���Z5;!�s���7�w���2=�rZ	3�*�R�2�hw�M:k���ɝ$&�=3�=6�&ۜeuV�w'����U�Tk]���-��n��V� >��
qJ o���A. ���G���a���T����)_��d��H����r�����/�A{I�T�ǐX�ϔ]��e���:�|��_���jY���Zk*c8|�a,j�h� �.ux_����mM��Q�[l	td� ��h�.����K���`�+�z��\{�a}����������@8��n=���X~�sC}�1�{E9r�"��AX� ��Rz9hB<񱈚���QC��0�K;(��c��vM�|������nk%��Ó��a���h������Y�je��E	�fW��Y�y�rh�z�b���@+�TӪ!�!?`���G�s4�]^�_�}o@���)����	��P�jL|��JZ�^:
<J������p���*�Ļ,C���10��Sf����� ^5s�S󍪓c:�/H�^ĝ�խ]��b�[�}��X�z5W���yN�S�A�D�Wh�,޿��x��ި����}r�^��0P��S���R&w�M�I��2M�]����1�1�&(}��os4���s]9��tl�׍sR#Ά� 1�Wv4�W����'p
�;�NL��( ��[5�Aǋ���|�˚%�R�~�N�^�Q���\�̓
q�g�!J�9��/��ř�7�+1=�LV�1�Z��Ė�y<��������r`9�lV+�̓*��7��PM�?Ψ����w��Z�r�/��g�8���/&�p�Y�i�M/=���t�7��r@�L�񳧘���R8��szd����I�<�^Ǳ�"#���A��cy�8)pH->��L���,�����
M���&o��	ЮF� ��6T��#�¹��l�cHmwJ���>оȌ���㧃����9�Pw��ɕy��Y��Wk阮��7J^JTD����ud�$q��	Tdelty�~���Y|�vxm�y}P�����5i��c<f�UJ�A�m�˒N�MG�`����ǉԨ��������In��ѻH���Ϳ��A�I�	D8���x�N��o����R��+ֺ*��IB3�#;G���e�E��ӱ�P�k�K�.���G>8ɻ��J`{����#ˇ~��k���9T��v8C�0LN�-ﺨ��^jH{v�P�m!�8�LJ&�/Y�jZ�1��m9g��2"��CG&�x!��>qJ�,�i������'O�#L�_"�g�}R{I�
%qJX�SP5u����ɳճ6��ũs#=L0J�P�-�rj	��� �_��[ڦ��z^���5%�'�(͏1�������4�䒳��n�nwH:q34��zД7w=��P<�>���u��0��
gZۜ�ym+��8If��
7?'}���I���9b�{D4�g^k�x~Y5���(���z���+�.�_�Z�W.Aۈ�|���x>>�+�rfɂ��%l�ص6�*&�Oީ��u����%�f���Ħ��;�q��\��ħ��W}O�b#%�N���fV/��q������n��"���P�'��cͼ�9(fs8:��ԝCq-�;��ۡ�x��I�F�<�r�A����eA�@R��S����=�z�_D��j���ޭ���/�l"�C�X(s�n%^�k�j+������ZDnJ��P�q�Ȳ|���@=��ܽ&>�=7gԳ-p;שb�[Z9ΰ�{�@۹l����Rfy�6���
?�j��'�B�!�6k�/e��<�ձ_��-Uꏦ���4Z�58榋-�Q�8B�^C�r�X$?�Ѯ&��ѽ��2B]��p"�qK��`D�c(����Ʌ!8p��p`��P>[]������s�L`��z�IHu�:JƿB!ن����֒2#�;�F����4� �o;�JH=n�B&}u4��A2ua|B_r=F�[O�R6jߙ%H���O1>�mU�i�Q>���~�p+|s%�j,m�@��\q�p���}S����7��P�D�~����Rb��M�4w[Q�K/���(�L��-��͒ѳ����SR�y��.�����-�=���[�X�T�ʋ��	B1k%���Ժ@���}	*��z%Դ�2���C�[�vi ��[3ъň�7���ar�d���P����F�iE��sӟ���%��f��T*�H���E�;C�*&�n���ʟ�q�MwE��9����)O�[�^>Ň � K�> ;�vd�����XXtv5�i��Ǜ�y'��B��5��{c�"��/	:)�
�MC���5h��7�A E^3��I1R��2`:6=c��]�G;��_���2J?�U$�r0��<�$�����K�y�/�B�`�b�j�\H����%)��e�̷��Kz�uڌ���F�m8@�8��oL�R������:� D���`n��a�Y�Mih�Z9��Ҙ��������]�F/� ���3�~�/3 +�W�6Z��+�?��6TJ��	(<,��s߸��q9�)kYF���^�m�zw����A"��캡��0F�x���1�>V��o�N /9)	��+YH65��JRm��hf��O�Ѭ&��\�@�c�q�Kd����H#.1=�	�mͽ�
�t����E[�q��m�q7��P�n�}C��\;3���L;�%I�B_�]�}U���`o�P<Df�Yd_�F�wv�J)e���	��`B��
��hqsŕ�=�X��s(�)�-w����@ �Կ3�g��X��Ffyt�s�V@:����-|�(�9���x��N'���5�a����ИdWNo���{�Y��GJ�U����+�u}颂�(���/oTP+���"�)��+�X��5&(�Q\�D���!��cU�,�K�=�{%V��=N,�2��\#����{�D�D�����'l�T�>��^�w��.�^��qG준�.���@`:kk���C��)���K@�\Z� s��uq�Z���ֿ���,�:�}X@�^ę��E�4w��UC�2��>%���G��g�O�wf=��I��O�\����/�D=����??����A>בF�ڸ+I�����R��wn�+gԸ�^�%N[H����2�{Ċ�~Ԗ/�iu��q��?�C-2���3p��kz���5�P0[o�s�s��9�L���Np*v�u���,���+����Lpß�9�+��p�sy8)��T�_�Q��dX�U���Q-_l�.u �7]kݒ��j�&M_ PP���K�1�O�P���Gj@-	��qß'@�e�4�4h5�p���C"����q ��Y���%��3ӳ��yѩ���=m�Q��'פk��6o�-m��H�6�]��f3:J�u�a�.��G�5u����%h(����o�
������"���L�p�e�=ZV��m�g$�&e(�Ǣ��T$R.��:���q�搢m��|�k�ut2�	ŷc�@TKzx�2��K+�:���3"8�%����>�,�N�H�Ѱe�l��\]�6ݰ�2�p}Y6�ù+8��_?՟�Hq�M��j?���ә��$�tUz>H*w�':��b(%�>����R�M�+�w�A$�_�4��� ��m�����wm���y��Զ��˕��?\;e����|)�Q8�Ј�?c?�(#&�j����q3k�|����|��]��C����PV�!g��I�y�����6�fT3�%����;��wr ů�<ݐ$�x9x��d���W�Z���ï!�GCH �0��"�b��B��ߪ���)�u�ե�F��@�Ȯ�D�H=L�PlI0�2�
0\�#Si����=�����蟍��XS�=�T�J��Vj�>��d� }zN:Q�")d0e �#�P����/EQ����4��7(��'hT�x��%Re�B@�]&A"B�`�i+*>�͞+W�U~����'�����GQ�����"�kJ :smh�p���t?��	)u;������b$��B��+Z1��P�~� A*ګ���K�^8H�1��/VL�i&����

ȑqikb�ȵ��?J�*[��.+]��tp��$��b��ڄ���V6�õ���E�6���[�����8w��/�Y���"A�8���y��W�
��b|I&0!7 Ŷ	��ܲ �LM7_��(��ブ��\�f�� ���|~2oP��?�y�K���ے�d����Ԅ���G8;$�z��8 ��Ԩ��U���/�3<����pt3P�w���W҉�'�b��(�َ����\p9��ͤ��辐�(ȣ�5�~������T�l�Q�!�Yt�4!hCv��Fo�h.(��*�[p#�i��}��h�߂���
5O�����֛lp��M.��6U��>Sg��(���,�+D	m�~qtի�C2w�8A��,��S�st��m�`_z�,	ق�l���?Zfǃ������V-`^y�jhY]Q�ۿ^&�HZ\��}�[aM�zYj_K 4�1=B�,��H�Ww���E�U��>�-��+%C�
��v�۪|�0�A�������S����	�3I�kn�(��̸��w��O��H�տ,$�37=�X]�@�.�L�̟J������/qW6�a�b*|-P�؋O����R���Un�+�D<�.�XT"�����i��6�#��V���hd���=�b<��=�lm�_FP�2���m��H	9j�2m-�b�l��K����M�ӏ���n����c_,H�o^�mV�h]f2�Wp9̩���L K�����aB���1�Օ*�A�X:�O9�h=���|>2�=�1��5P�O#�M�~�V_$�� ];L��{m����4o�h
��W����֕jG�_��v;Y0{ET�V���Bp�i�6.t�����}� �[e�$U�zB����W��$T0�� ���2��Y�_Җ�@kW�h{�n�e)/RM%+)X^���L�qPP��Ǳ{�)K:!+��&Ǹ`�`��T�HG�����]K�h��[(_�*��=7���x<p$o��qU����V���a@�NKh�]��`�G�z|x�5pp�M'��r�0R�g���+�㸳�ik��d��6�SD`�;���!D�X��$�$2�)�A��wݚ�粱���m7�gg�B�z�ڹ��D=Y�.B���Ԍ���%w���&Y�L������M��o@�"����E�$�nvt	�l�����C"�y �u���RA��,�Y�~#�1C��5�M��C��&~��"dg�QQV��H��^tUM�"Y��6+L�w�g�d��A����YW��ǀ	6��f$n0ǳM�����p#����[$��p�Z�B?{������駭�~W�����x ꒪��,\0&Slh�ӑ���F��ۚ��`�>r�|�ڼ���)#��s`!;���0�WЄ?7�.��_�k ����yL[�Brcc=��ϥ����םJ��t�ؖ�@�n#c�w09���2��b��!�u���[��y�6��%KT�;���&�u�?�XkcD�V�Q��yRxe
���:�n e�'�&J��ʈ�O��xܼ �9�G�-���IT�2�=��W�߈cmn�gY�.�yi��@S����tn|?���~����:6S)����
�(׬^܃���}S��*�X���aϑ�f�,)�����r�h�4�Ճ8i^��"�eJ���3�1:r�m���T�~�(��ܪ^�3r��Sx����owA�<%��p�~~2+��YqqOw�D��b��M�p!���qZ��4��qo���V:N�-PmlU_�'t�I�ꠎ�����ܙ�z!drz>5��Atɿ�!�=kG.�:��<�� S>q��M���u��0Ytyx�Lu�y|̔P�^߼c#V���!\�Au�Ou�R�j�]�
Ԏv��>V�-&0�E�N��	�>�!��a���,4Y­s�z~<�t?�V��
m��/�����$�I�u�l�#鵂7����,�D�K�rj�i�ig_	��b��Y5e8��RLQֱ�$�? �b�@�=�j
b�j`v;��-�2/����m�\ތosv���Y�'h���G^�f�܋���D��Z$"�<�Se�6��Ӣ�����;�Q����r�T���ʽt��F��aCM�fU{\l�U��#�3��v��E���W��~��ܪ�w�>�����IM^��{c"JX]8}�A�y��U���U-k���q�W��E@	�'�`ӯ��s�X���
<���w��]�T��sj1�Y�J&y5��lȞ{�(݈�q��'�Y_��acq����n{��PT=;;��d���d��y��S��j���F�|�j���mJ�Kt��F& Yq��`�t��Wѳ<0t���R��Ԣ�g��k,a� ��z��d�6��g��Fx�ĉ�^Br"G��6�f��6ᛍG���rG�bO��N{2�a ��5
���y�}�yl�%n��P=�Vҋ댹��d�����q3<�&
Z�[)a�<�P��1����.v�bӛaV� ��,�Um"�ޫ@������8�%>�DW�2���`�*�?��؞`]���L���[ϋ���A�2����O�|�f�U����}Wt2��Zi��*��{dYi�e�!��x�?��i�e=�H6Ҭ��вM㬕q�����g'?BR�H�
��"3~Ͽ�SM(-qO9;w�hl�"�C�}tR%��e׹�ς���o�連�!=�	�����d$W�ǩ�xS��@"�Z �b�N%�I!Y��K���G{��~��m;N	Q[���(�w��`
ې/��f~�ķ� �^�u�Ǔ�{���c)��ټ�;lT'{��9N���U��\8(����$��I����\(څ�[1�Z��P��+�6�N�P{�ڮ�]#����~rS�����v���/r6���m_ۑ�Cd��z��ȀO^~q��~���p�r=,���t-3����״(�ۥ��:�_�kE���G��857�i��?;�k5����2�����W�Dm�?5�P����I�@%X*�Ԁ�X7�m'��&͋ց]�D��wU�'�6wY^s	D��9�Q��� �����O�}���Kr�#�����0��Y'��<l�M����8��S�s��0춱�P��;8�:�iAm�S�؊"l�N�`5�7#2�+��Q��|�*7?x�ELϨ���S��I�3�#w>4���R	�[�
���w�	1n���r��)��V��j��h\|NE����RḰ�#��3͇�6 N�%�U^�T셴�~hv1�U=����%o���U������T2�Z�{h��5��p��^(����q�씳��<q � ���nGݣ�쫃Vi@8�XS�#9%��_+f��|Y7 ��h?^�sx�Zǅ�8EFB��ɂ&�)v�[�E�����{��+�R�9.Z{�K�k��2��Ս(!ڂ�����0p1�5��i>���K�D=,;t=QuLJt�3mx��%8���vT������2}"��Z�()�� .��
Q�K.�g�~ �!�^3��jbkH�������M;ǗS�K�6W[�T�1�I��J��1��C�tv���p�h����>�K�u4Ԇ������D��Ix=��F�@o�5+b*S���;���Z����F��1��ɚpG�����X7~��2����bv�ta-�^[�!md���v����� @��V��6m�<i�^���bȟh�E�S�m����a�(��;2�1�8�/��ٻ�[V��Z���9r��QT��7�.���/�r�-���x4�AE�:գ�)����ug	!DW�ڭ#u�?�����Q�ۋ"F�R'x�"�'��K��9%Z�E�=��N�׵rR��2�3�?����&K*	���IW�߈���w+��=�����.�34�j}�.�8�����ue���yM��&�bS�?�r7=ζb�����z��݃H�Q�:(���#���k=��L2�Y�Y'+VL�@6��(?҆h	��.o���Q,h�	ksΞ|�|�5�
A�z�ɼ��*P�f�l\do�?�-��	�C@ Rd��&������qɇ�ϫ�_D�� �>�x>��h#�9���s?^&��s]G�p�*"l�h���͔lОx����W$�ҙIkĎ
t��\����}������ R��`@?OyS7!��=TwA�Gk�î"�,��ش�p�k8@�&Н�p{�t�b#�?F-��Ԍ���2_"J�m�y�!��׹�
�;_Jn�n�릀9JT�nk��>1����${��g�o�b«�iV���f�2��nb��\�$��c-���ష�V3�f�J��W�H�]H12O��,O�bk��.80k��е�P�� �G�Y�.��}S���dw5��f���g�5�Y�F��rߍʴ�B��gi>����$I��1�R�|�6�>Tn)���r���_�*M����ѽ�A�P�l�S��e*��-��101�'#b����:�� �2p�H��=a2l�-Ԛʼ����*XB�G�B[6و�ؗ~�����U몉��\M$��R��qC!�w0��_~w2��Q�2�>�"��q�xŖ^*Ϭ{^�!�}Hp��}�X���J�p�������B����D��o���MV��������+��TEHqZr�6�5�$u��1s��,V�3j����;IF�YPC���Gľ�c{`���߽���%�e��_1�r]��Ō@v��?bx�-�6l�&��d���H6<FX��}�G�{X%)܇�T��x`�?��i�(�b��A�	��|���ܰ6�`�S�����=�Jj1j�۽�珱���z#��; �%֣�'��LaQL�Ş�o�EA���cTf��r���0g��I�~�Y[�b
n��Q���S�5*a�I�C��|��5N�]=�кW�z��`<j���F���_�.��YQ�$|A5�1�brDu�Iy��N�%�k�'��`�u{r�W�v��Y�8�2Ǳ��0e���d�*�?>������b��-&4Y
w32`:�ϳ��gd�O��8⋱=�3Q�D�|��szq���r��r(�=��=�rN�mX>_��heD���N=��\~����v��D��<��.z~	��i�&�NN�Ku�)>��sz���9��c�b�*��[�Tn$�Y~�w}�9?Yu��Ě�ܟ��g�p�pc�}k �ے�z��]*��������1A/*r͋�Kn�Xk�d��H6���3���*Ϝ�q��Q'B2��N�����bx;8�4y$���>��夋�W��X���gv�,	�6:m�����~�؇�+�].t7U��6g�nt��2����ꧽ٣���	��D�Ӥ�2�I�����`E;�"�D� r5e��c�[wF"o�O��ʉ���Y�2-�Q�?�t��j�%d�B1o�uӰJ����eJ	��<۲�)Ӈ\PP�#�s�d<��!��l3�&��g�{j9}�H0�Z�8By��oF�DC	�+�j���e���3t�>�'�$6�����|q�\��=�߶z*��p��+�����~䴜.$u� �%����$�u�p��*r��n�DJ3�2��-&�]�����/��k���ғ��C��n�(�j�6R�a�8���I�R�J@|�S�� nT���ɟzYd'��	�U�[d����㼍�S�F���_KIldTffW�����,|x�����L�""�il��Ѥ�w5Z<>̖�uj�ǽ	w���]^����-e<����1(�ڢC�N��l��S���N�W#TB��_D�H�aF�>e��yJ�l�A�~FL��D�H�謆{C�iы��u�7ɣ�Ud�� ��q
�Dc�ޔ|U�;R;`�)\0�"J�H�*�E}2o"�\����!qf��A� y��6�H3�*�jʭ�����;�V?g�i���+�eFz�������VG5@�TRs7ܗ�Wnw�C�J����Fr���[���o�oTh���5Q.5.���R5�Ƶ?J���fe�Z�͉:D
�.i	*�z��.��#��`���d��5�����i����)*�q	x�7;��"9!���v�Ib*:|G�j$�hV��8ԧ�M�`=iaV��J���%��gc�n����ʍ��$�6@נ�{D�f��3~���r}$����-��UE�T�Rn4AEBCu5�p	�G���� +˱�[�]�I�r݉ļYtT�ĳ��b����KZ-���gp�,�p�;`�r)ZDf?aǁ���/B����3���I�Q��*������*��wf�5����6zf���$a'���-z7��\ñ!0��*j,�U�*��FH��_�TW��Îk��\rnI��t2Ne�
��s��P:��t���<����,�59Q;X%M�3�`�&GY�l�7�mZ�&�
�l?ۇ\�H�ca8�vw��"���^e�ʣ�	f������j�i� �����+�5+�%�Y֖��>����0Vz`<������*k2��z���'H��0�3�y�=��/!gT�0|mŜeW�����ϣ�3)��0OtH�@��G�޹�&/�u��N�+)�.�x��=v�#�,Q��J�p�HQ]=���6�H�ڗJ�����w�?x�����dK��4۱��y�b��M��
Fc���a����J\`�[g /�,�m�޼�4ƥ��L�(Q���WFkqr��:[zcï�x�\vu�Akv ��@�+� �(x��V@)p�|Ԓ�9�]�|B�N�F�O��M�I�ٌ*uP�L}��:�	n��1�Rd��X2�c���ZwL�\Ӥ�BPZ�S�֕�j~]����b��38�+�`�v�d�J�xpL#:K��� e;�AwEW�-�K�nY�׊l��Sى��;�;I|��ږb�� ��t=��N�g�I��'�P�?�/J�z		���֣st��k�(�d���V�����Y��D2�8����f��o��*Hw2�nY�|��A�����g��ηP�����I���̡�=�=�C	�43Đi�y8R���G�W
�>��|��ے���;e�nV=c��-�Ǩ���*��-O<O$y��!W*�o��8��0��
�Q9l�ki�['�'��������[scǦ�ɛ0��¼��gJ����y����yy�m6�q?������T���V�Zi��I��C;A� 3�}O@`=��g��N&�*�i�\<��P0��x��R!S�]ߣ�o8�@���C{۶���?�:��CE�����.�h���ZC�����T�J�AlmoJ���j�h�T��E��F~� I����8	Í�ۺ�촃y�)7�����.��AKۍ��r�ō*��*~�����닽8I��Z�N��v��)�=$���P�p��v^�t�Ad�N�S>��j]�t����#fk�1b$���g~S 2ޢ2�B��U�X�b:��7&�ܗ�����y�`#R�/���8�=�俴N�^�>G���c9�6�:��^l��b��t
���Y�>7�gp#a�a�87�'�}���s#��}�����s]ds7�T@�wMâ�_܎[��mQ�H�'�e���������OM]T�fyA�z���Fq�������z�9g��gN!tz_��`�W�ofɂ�Ȁ����Nt�Zqc��7f��WV��d�4RjZ��T#��ѵ5�#��DOj^�"��Gw�WNQK�X�z�0c�&��RAč`c��v�T ��5ry�i��^=9��Q�x�|�qGi_I��ݶ���:�Cw���`�W�5U��V�ae�K����~��ϛ�GJ�c�ջ�צ�c��!+A;��R��<����!������^��"��<�� ���%�S��MS��3f�6S��L�6��ʆJH�f;}�C^�"�4���.�x�_z0ph�mL �<����C
�v�χ�i{j��n.�h�3��ӯ���	q�a:�H�-��h������	��v�1�[��C�j�N���L��Wp:J�c��+��YM!p B�J��k���T~'�{��Ԟ�fW?v�f�^E6@�ϸW�&��T�$j��@Ԙi�7x[��i9�p�o�
���wY�O��n�]���|.���w���
2RO�m����{�M�1T����k[��R�X,��nvc����u:*(@�HnW�3Ff��k=x�c5X���˭�KO]���]��BY�^O{mh� �)�T��"k.�m���[�k^ 's�6
�)P���w�-�俀�8;˛�\:-�A��
����Jo�c�����3�x|Бߪ���&�ƩzKu����T��4Ճ����/����:!��� Bg���09�D$nK/d�,�p�e��H�M4S�)��yl�-���٣���"GYÂR4��4�֔x�@�b=�r�16�7,i� %���(�4!��,>zr���#��tϱƮ(���.��n�)�����"�7��L/V�\�fݤ�����@�T�z�=�l5�f��b�Ot �*{��S��Y��eY��]���F���i���G9�������ⲨB��8|$�ȻYD%^�?������N0��!�=���JFzِ[��'�ǳt�^i(Zz&+_�W�����=
q��	�Ʋ=��f������ �Ν|��x�����%I��7N�����a�崮�.�;O�~S�@W�� ��7\�>&�د��xi�E�8�7��P){�9Q��K����Ҁ:����Má@�8H���D`�G�'���`h9�����U뻽�ZTeEoK������,��"ד��Gp�x��P�H�'EmH�.�舟��״�m��W4�q�X~m���NA��\kt���mJ�0 }��(�Fj�if�LƤ|{׫e�CT��26�VX]g3wC6Q��\�`��`�������=X�#XH/�+�`3o$����З+x�@� lUȻ�7r]�#��#e.�D$�
�s�@�:�d�"��򛚑B�)N5��5��>���,w)�Β*�¦H'��$S�!��xJ�c]�2;Ud���r�E�ۘme��oȳM���p�G�P��?A���n�5����q��k6(=��0\���jBt�v5}u6�����v��f�A�0�:K�����ó\
�@�Dی+��T:��8f/cX9�.���$0��_��j&���N�D�s<����	k4��>n� ��!IA$Sw���Gm7�C��q��?s�j�?�Og縝�<�H�{���-���n�����qH1W�6����-!֧������'�0g4`MT��
�҇���C#3ʨ�+	n�q������#���i<��/��y�7��{���L�"���m�#V�����I��W����T�d8��L���W�-�8PkG�}������J��6>Vg� �e�:�ʠ�1�7Qr+�`P��;M^�_��tA܅v�%�
�����������	b�Spj?���x	*.I�K5����1��fL�����DU�yl�hn�Z�QJ��@ε�N���f8.��:���M(�1ы�)i�7�"�������UZ��x�k`_�2�y�L�eMg|N��#&���S��*������>#+�n�uڀ��"o��f!�j�B6�}=���煱����(�~B���xB��&�4Ԧ�+���>{o��]%�T\9�+����@XR2�"��u�Vv,1���;�e�t5[��}��H-�.����t 1������>��2�<��ܜ��OU���!e�<?."�!OE������%�N�Sudp�� \e�YD�2E��sg�ѧl^��T�؊?���t	�����74a6��,�Qa�5�|a���A�L�������" "�"E�.�$52�	��$���&c|�'��=���{g��`\h(�b����+�r��fnogSrg�E�Ҙ�'�g��@V�T��@rG#��2?�W
��̎�}N(;@�*�VC�������I�սx���<@�Ǉ�6	n�&��N���8 h�$d��%~�z�&��;�|��#)T��#&d���%���t$XX$����mg��p�}Q����d�����ʒp8�E
��ˡ�2VN7�"oI����Z5�3̸6i��6B�شZ/��R@jT?h����~�8m�Ol��)�A�$C��y�,����#�`2�e��Smq���\��bx��1���9s��������"�f5�V�T�T�z���ɉ-R=;�	�3/���)э#�e74�2��$�E�u��$g��5����q.��~Xt��7'�3�BѲ�\��mC�1�h���Cw�[��n�D��PI�:l����:oShɗ���?p1��=x�z�̈́Z�ş<c�P�/Ĳ�� �\�ҩ��9�\|o'�N��������Y$�B��o�sx��
��m�'�;ΰ�3��A�pUy�1I�!ߎ��4뗰�^|����^���;p��$���2�����7@O����_�p��Kx�Vyh���b�]�ꉻKU*i�$w�4�i�;S�ӎa;kh����L��@�D�4�A?qq�
���� G��	�Y�w�B��i_F;�@L9]y��+����X�r!���SA\�B�®>�[��E�����j͆uכB��-��TQ��BEL^�����|5*��d�Q?��开ō�Z�c�"�	N��D�b�8(
����H�Y-�Ψ�e�f5[w�K�N�rd���� P���;�]��Ⲁ� ��q r����PZ�X*na:&o�tN�����O�:�xA�Q�S�B^H�Lc�94g4g r�9R*#|.��y�*0Lr�`Tf��?�����c���zih���q	=�9O�vdb;�:0����H����d�!^��ɓ����<tYc��9AĭX]V�D��NT��k��q i�Fܒ�_<c�L'w�{F�5����ܰ�g��=�����l�R廋~��W��yѠB�c���R�/��|���{�kې��U: S*M����8�C�����c�7��p?�&o9�h��+�0϶Y�`�f7\�q�B�@�/Hb�yǺ��$*�ʔ�[*QQ2�;�G�w��N��C�W6��DS����LK��+2���<Ղ�ޅ��!S��H���eA�P�HDů:Ï�d������A��#}�" �Z&��@G
��������q_"��c�j73ˡa;���sZJ�YD���Co!��`
t�QX��~��Z9� ���@?�x���{�#HaFQ�ͩ��v�Tƃ���m(�Uniؙ	cs/�7��/�ס^�mSI.L������u�>���Tx��3��1(s%E��}>�ѡG5N�i
�ƭ�DwY��}��j����;P�s&�h�!���+e�S7�@�'g�iAj~���ssW�*�.{�}��%�e���b��N[�hd��30�/��@^�7qZg�k�n�<�]Cvtw[��ԇ��hP�'�����B�8"՛��opw�؅���;���W?0������d:�� p[_����"���HTzTxn��؆�E2�����'�J�~VS]`��6��20Љ'�};A���Gf�u�ս1�R�N�Xi��x<�R����n�@.�݈k
��Һ&��=�h?�À$����\ޢ�_@�S�{ۘ����2xS\Dנ��7��[jMb"�n����V�i�[������L?C:��Yd����*���Χ��K*���oV71�eo��I���$^��{�s�[���L�x�,��
+j�V0��I&k�q�!!�j��ҥ$�~~�R���e���ĭ��(Ke�oH��y-�����4J) t�S��^�E]�8� ���8T�.��&h��ǭ���?�6'�C�Fźm:5�5�����[��8�pwhf��^�`_���ś,�]�(��D���x%�qN�@>��O�tm�7ON����;��A�� w��UL��R#'��S��l�>�kߓ�>����ݜkR]1�39]Hv^����	 ɵT��(����:?s����
ޑXV�'~'���� 샣�*D^}������c��/�)E�O����n�#�����h�=��Y?fW� ������]���i^lh�W���>���Hn;�r�Ŕ��3(�>q�����o�4s��+�Y{�ݱ��ݖ��	��P�c�J\�1a��B��'v-��bW�|�R�=<���,�9�'�Y}�������`Y�J����P[T4�E�{�tK�����Y�IA�}���,v���N(�z���W��o��m���>�-��\��^�H"�~ʲ�����!=�/��u?�,���.tM~�ⅼ�������K^�!l�Rg�>�����jZ6N�V�܊�"�^h;��^4�_���>� ��W뒼�j�S����,��vΕK���R�RMMV��L�X��Wu؜����������j�&�J��%���5��+�nK�h�bI���.ޓ쟿���qP�k#�M у�~%ސ!D.}����	yTiu�?��>lKp�'#?r�(mX��r)I';W���w�h�C1��vC�r�{�mA�U9�L����ۭ|d����*�]�Ɔ����#vE�=��7 � ٍp��J��)a������RS�jy����56�� ��&�K� ؐ��?���Uү���[�Z\�@��|�R�sWDb"Z�f�d�L�rI���G�f��<}QD�,�H�_SfT �@׀��н7{Z=�8�>���?` *�ۑ���o��94��W�Xl4((�:��YO8�.\@�ną9���;�~>�iP��<S̛�S!Ż��f]����ߚ�����;�.	�\�L��rk��UMF��.8F�`�����D�<C���UClb��>�����<������g���U&d֩:���i��w$��cҠ�׈�N�~���F
Zm�<�-�#l��Z񦑜rP^�3��գ�l�{�z�-G����a�š�ie�#�[6G�]
K�������L�/��]���l�< +�{�s�<��K��_��{�Y��D�5��3\��) �����,����l
����[������	�S]6�����Li:�)��ԈS�=I�g��k(�@��6���'�Oa��F�X̙/�c�O�,oɀ{�^K�2��d���C��٨ @Tʡ���Q^vDff�y��t�ޤ@K������q ��n��yE�6�;��F��h��yՌX���o�zZ�TS�@�:�#T�u�G'�?���� 2�@�Ex!Pj�Wq[{�%RDpxJpe�m�?�8�#$<�'�� 8�0&�cGQ�lk$[�?�������*M����x�l[o������.g��L������%b&
�'�N3����2_M٫�����R!������Xr�F�$�n�i�s��??m/N�"ǪL�Ě��Te~��-����ꭔB8	Hzo�^�ƫò�����=���@�S� ���f�Fq����@����V���2go�Vp;�c�ȭ������VŇD�ے[�]u�T<����zhM(�3�*����4��.q�N�L"@��U%���������nT���8�+�47�wV�h�Y�i�6Z�[���C��Ű�Q���0�	�ETjzC�h�/%S��V��X�;��W��[���n���/(RN@���
����ǝ��(�s��Q����je�W�x7OY^�c��*���_�U#s��1�����y]��*�H�80{��i�]�%l%�m��!"��J����|ϏI��V]ȉ{)�T}��u�8�l�"�a!���!��l���%I���J��?�yeLl�g�O�̅m�20���3k�Զ��{�#K\�s�Ȉ^��E$����ƕ@Z�G`8�C!�U%�垢������̾�-�I����0ԶJC�&�Y���ֈ}L�6�ο~�sƒ���J�����E����%� �,�wU��?�R�F@ҳ�~��z.a��[a��Vc����`v��0!����W�������j��ڦ:K��T�Jh�W����Q�_���$�`� ۷F��b�噋I����.���g���R�F�5�#K���!�i�Ld����B�������[���&��Ӝ|J�ug�rjS�oh�*,���C�S�=�ОMGz�3J1q�WPQ�ɐ?.X�G���s���w�_L��m}�+�����Z��&�j�p5������w/V��zn���$Hp��J[�*t�G&��1��=���1{�/��l�jz]��E_8 zh�ͱI�a��:��7���ż6�㨟+��*!M$�t�dꑮ?�HF��u!�.U�j��(1�ZЁ %��c�'yȰ���b�r�RQH��$4	����;$�n��o�P�H,lWP9��8�`8ka��=�A�ZX�&n1�O�6O���,�6'�a,\�{%x�(i<U._]-���|2hB�����a�P�~0�ϰ����*G��W��gb ku�FѺ�"G��uw�Ѓ_+�� ���ړ3^^P�Z�<	���w.���%����- �ુ�]>E���i��Z�Dk�n�%��-|��-~#��d���M��r��cX���Ęx9��@HjѸ�y�8�#�9���7Ҽ����޳O�,�L��$|�����>��(<�zG>�/�����IH�+AX�� ��A��r�V�n������ō�\ŗ�#p��	˜�Ѓ��p��t�:C�I��n���H�$ݟJ�!���)����s�;�jy_�29\ME��ͣ1K��T�"�ޮ������̪S�BM��r:ݪ��H0:2��и
c�X��de��X��.�����̊�k��ځQ�ht6>Vs���l�� ���K���W��	���A��s�nY!v �??6	/|U�f]h���Hk�~xhX�/v�{���xh�x�C�����L���ju,3��1�XR��wR�bY�����3�k��5_>�KD<�d]XX�-pZ@<�iOQ�c�/fkX���Ocf���v������n��#ӣ���w��Tw�g;hTM[��l��vcͱ�c]����y��`�D�����)-�G�M�D��ZPJ��BG/�~�c�G&�
��V���ֳ���d|6b��g���w\_����Ն��z���W��a���J�(����e�Ǚ�Y��M|?)-���m�k�>q�tr:t��t��e7x)�>��X�:����1���1�_��j��0�	���_��%����6��g���˚|mH>�P"[M!j������Zb�*�C�oA9(���s�)�g�^D�	bn����}�ث7Y�g��.9bDP�p؊��7־g��]�֘���0X�\9ҵ!h4F�������$���s���ݢ�t>m��iA�D�?ݹ�nCʯC� �Ox�\r����y�x$��ܮ�{A%+�MX���Ȑ�<�*7��|����ˀLg�$�U��c�������%�{if�y�T�Җ��?��7����eQ���7�� PS�=�Yx�Q��ڙs�$P(
�Cjo�9]4�~����A�� �N���H_K��s^@N��f�zi'�1�c�1|�� ���9�ILߙ'l��Z�@x�Y�l�G0&��_=�m̮K¦áj����n@+�s�g����5�x��xn��!pr<����A���$���pPq�1~_E�:�����PR�$�$��$�6m8��/�����èc�ɧB����K��Фm����y�u�@b*��C =&�Aɡ݉�N�ؗ.r|�eoQ��g�r����N�yyG��bh }v�H+���(��X.M|�=x��
:�+`"���!0ΰ�:��e�/����^�"��j�ޫ���c0��э�>Jͤ�oa�eW�0�x��˃�t��h�[����#c��D�gűqt����Z�n����b�4�nv�Y�8�q�[E�P]r��������z1�W�p�[�c�V$�߂=O�h�ki\��~Q`�|��m��%vD�����i;0�篥����p�m�;�;a�����sKF@4�c�H;M"���]���%M�kA�=f�d\��|����s�P_�S�x0�FgMIx��v)��~L|�Y�V3ZD����C�M���������9�L�[�z�h�#�ێP��9��4��J��t�����Zj���o����C6:�djr�v�A����G-`q���������2d�F�'o�x(�3�њ>�c��pi�ga���y3j1�1�m�p�`���ho"�e9c��	�S)eh:�C�\0	3�^*`�c O��ȨL:=�%k�^7�0T�e�M��[�$$��ܗ�iQ�T�to���u�<��h/h,]�/��J�c�{i��S����.	��BM�ݣ�{��<�*)i'=��1��N����(�����mY@1A����aPƴU��tC��������%'@��eZ�ݬ!-E�̝5�S|�KU�cǰCj��ݑ�=[��HV?����&���qP��p4|��f$���D������kNWhcӸA-\��۷�����LIp��l���y�˅�gƎ�%$ŭ�|fq�o�?�$s�����Z1�J`.�hN�4
�;�W�q[�~���TT+�&�#K��cz&r��f��vo��zv9 Ŵ|�Ҹnk���4����z�Dv{�ii4bNYJ��ټ�4�)1���}���݃�iiΒ�FG����v�U�@��z�4�\LC���|��mvmo	�����)�J����my�������ضx�~�u��q�ӆ�^�rBG�Z�[��P�,�{H�|5VɨyX?hZX���#�VT^�Q��\�0İ���Iμ�|�
��S��"�M�%L(��T�2��_�mz:�C߉��k��ָ�A&���ip3�L\�Ζ8 �PlA�,։�d@�B ������gz���V�Е��qlt
$��;T�Y?�)<�����	��I�*��d|���T\�znZ������o0v� ���G�����0��m@�� ?��O#{D����P��j� ݦ����?9q3Ȋ~�tWD>=��*A{.�� y��mro�1 +K����tu鉚
�Jp��jҙ��Ą|ċxه�Z�g(�X�j��;�V��y��Sa�����pWSO�#��~���e�h���bK�������{��X�a��j�	_��&MA����N9��!�&/a��� �zJ;�"%o����i����5�3(�����a�c��P��(]8U���._����(j���ᝂ]FO�E�:�Ѻy-Z�
��)״P��O`%�^@�>A�ֳcy �toa��}���H��^�N�!�<U�^�#�H�v�U�:䁢O:�[ow$8�B��� �ؔA���!ݟ��+��r]�0,�#V��h��d�dٕT�W_=S� rS �fU�b��˞�AI�kb�Gz[�z��ї�W��W��H1{�pxQn�eU?"vz�۵@%�Yr���MI��nk~Q1p����ӥ��!(D�[��(w��)`|�"[ٯ8O~2�����<��~i�^��+�<L<��[�s��7�����d���P���d~:��o����]j�^�V�Pxv�'O�}˳{N���m���B���*��E3�m{dUQlk��[)�'�z"~��`�S��j�h�y�Eb�.W���&>��A�e<S&F=�F���gu����hiu� k��������T�Z�і|��=l��W4��84�xU�t�)��1��ʙ��Y[�E7iK��Hy�4k�l��}(`T髞6����zE��t����d��VF�H\�L�>��T3�Ψ�:����M��K�������c�-j����X	e$ <���|��Xg���
p��`���PԊˁ�w��Jґ8�!��h6��eY�`�/Z���H=�|HH#�(�|��q�9�z�^vޢ3���"�o��e�9�uW��'3?�
̵6*fK%�w�(�D�A���L#Hk���N���l�#��`��"E|���ٹE.�2�s�ڴ���	��W[A�S��t �=#�B=�2b�BU���.Y�oz�GU&u|�U�������o9X�ٶ0��b$���A@ql�I���>��r�� V�\�jM�D-�>Ǥ=�u'�H$��&�����]u�w������.b�����Į���9+�����X.��2q	���//�|t��gt'�M%J&�!9�VY6+L�	Pw.���e������ܧ�^��N��.I/��#�m��6<(2��<&qV��"�/A@u��,ٽ��?�PF�ԗ�K�]���+�	D�C����bԣ��
~�@$'��M�H�C��H�Qrw�	D̪������G>N2�G��'�LZ�xQ.r�
���v��Mo�4 Z��,9P*KFPc�o.���E^���J��jm�m��l^|M�*@���\M{����ŷ�ck��O��!o����4v��X����
�<a���������oASg��po�I7ݑ0��S+���t��lnc����0$?Eqq��R5T끺�R�	�n�����KB�,o�HV��-&��[H���enz@ p;��:�GCx�p�Ï'�N@�{h�"u����\4^.ӏ��$���Wo��JFk�#7�c��_\%����3F�� y���xI���1#��>���V�V?�a/�h�v] ���?Ѕn��Lk�S D_aa�E�Z�z"�.�M_9Z�)=T���ìˀ�P��F�f�I�0�����	����bթ(7�;�g-�SԵe�R�����J'����B�Q��b?sZ��KcRZ��1��<$���S}�^ 7l�^21�-"r��F�>u$�Q� `2�Ӳ�Y���|��9�W�;o�2NG�����\����φ^�m�x��V8�s�P����ԭ=>� �7�>�}�ϹXV�H��O���~�4/}�`a�\���q
- �������.8ҿ���[��b��VD�&�M��m���H�aR$$�u�H�������p�g�B��q=R��C�o�X�̣2�@�����0Z?�Z@�fmukWM�����V�;N���QO ��
�{��U߳d�c���� �]dO|W������(�h������6��i�RX	m��)������P���'���"
�w�]<���}������U�:��:�tS�|`=�B��,H\]�k��堛{BҒ˛be�f��sZ�
x[7�{	YJ�(�j�f��F�v��p�}.�ɯa�)Ɓ+�t�P�w�zk,9��2\1x+���M������8R$8�C��1�o�k����Z�_�s��NՀ�(��}�A��OJ�]ڶ�S�dn��pZQI7n.Xw���0X}ts}�����\A�Pn��W�j�;��hg& _�W��f�Y����q�m$&Ɛ��{0�4Ƞ�(D�j-��"���툀���:П��_��������o��=!@V���'i�<D���I�%�\>����rc����@��b���5�bTp��"�d���j��ir��qԃ<����.�c��9fp�1]p�%er3*��A9*��]�,�H19����:��N��Țd�虨�&|�v����D�?z7�b�7߶(;}�5���6���,C��X�!�IA8vd��4���-�	P��s[\���k�=D��{�>#H}��T�E�ۧ�RO�c�3��F�3�ZC��	��Z����xz�x���?�G�$���x���{մÔ6[����O(/O�Z֍����V�ƪvY�#�a9��(Eע@7���
u�����ݝh%	��1M��І���wb�<L7-�>�`*|uh�q�wn���S�)�C;��mKC�&/c��	[i�+ėi��!�Ɓ:0n �8��-1�JrK�ntWG���kz���%��x�]K&��)�XX`�e���Eˍ�l��tȮ�>RngZ�z yZ��e�u�=�P�?U%��zf� ]�|�<��'��ۅ�,�8w@a��2ØEU(]�I4M�{�Eڨ�@b6a i�)-/���}ǂ �w$�w�����p���8l�7n���Fvͻ�����[���^W��"̃�j,�2�l�z1���l8b�N�F�#u��p�R�d�E��ֳ�"1lj��^-v���3�#}l'8��B��[�÷#j%�s�@���ވ��I�՟�	b�|M?K2ku1��U��i��sEê�;;ӄ_�:/3�L����R�����5 �4��⋍)YԐ�
F�]|3޸�~�+�$�����b�?oYy�'{D�.{ r	�"Ѹ�ٺX9��Ĵq��� �9`�NM'J3.�/5P J W�Np�!�cƓQ,�ľ���G?�g����t�9�{��Y�8����ԝ�K�T�_�H�t62,*n���ԭ-�r�=|�Ǎ]�Ⱦ�-/,�ŝ�:��ic=Γ:h��U=�K�Y�M0�C��$e���7[W&���ƞx�����/v���_�n�m�Vͧ�t�J~B��dl���1�g|��7�(���N���ͧ:Ӡ� �qb{�����ށ=b7=�Dܵ :��Q��G���$*KHH�������|�X
ۋԙ�$������P]ޥ��h�RTj�c	�϶�1�0�+�f�e��I�$]*]'��?��PA�2i�/�\�h}**�=m��OwdOz+�������o�VpZ��k��4#�Z���nGxs�z�q67�.v���Sf�L��{�EzRw<����=�S�|������u��z�����:�/�D��~bzY"��t�m�V��a����`(K��/������o3�M�f�q,y���=LNZCi��)�z%?.zGm�x�V�9\ԉ����h��7n�#L��{�B��L]�̫2,8O��7���d�3{��A�����S�z��]Cd=y�]2R��]�Ɍ�`���б���8�ʋP��bH�pnL��~G��p�25.�T>�ąNa$�Q�[ept!�Z�؋C��N�
��9rG�6·�	�q��3��Su1�ŵT$�q��BR��ʓ�P[�M����ܳ�S��Lԗ�8���ٌ4�QU��.����X��X��������j�b�+�yY�ZΏ�����[o�-��n��N~�ɝ�w�CT	�`����������Ā�@Ԋe�϶`�d1�HW�Y�"H�}�SOi�r*m�99#��R�Ɗ�̿�l�3S���S���7�^�-���"�>�Y��#F�4(�d-u��㹠���8���?EX��r�q.���il�����m֓�Q^�>�7��-�s|�+��F��+K�!��(6Q�SW�E]�����R�gj>RK�L��n�2����^̖jf�M�����\k���C�.�D����iQq���S��rPI���M%���i?����f��Gӝe�\ټz{_� A?�h�����������<ޏ
�H�B/Ә�+��B
�("��Ydl�c�<�W*H��� ���4��y�衕/ҧo�~�#��
��)�KSf���ʉ@�t��V�/hH��:����[H��'@D&�,�H��r"8`mo�E�����tl��ӟ1D�;
˃@|Ȁl�8� �T�.�B���C���!f'�	%����w*J���޿j�EOCM��Y!G�7 ���ux�nYr���ߢT��&�J¯��+J��\yHW[�O�m��N�R���c8�Pe�{m�9.a�@j�O�k#쫡��{��U���$63+�!~5p�}�\�	�h����`#	덤��io������,Bt�=Y�`�a$V�9�������D��Ţ��?��Z��V������4�ȍ��r�{3��	7��=�5�m�l࿻t���Q'���n���R�����`�H>l�'�9�2���N�R{@�
1�����	�gi+���J7��f�A�_�J��Fj��[ge_�"C �c��@۫m7����IZ;}��З�,��!Vi�R;f73�^����z!ƺ�6���-�FD7�1��&�%����A$�gM�P�E	����� ��(� P���R��zbV�O8�bN��Oj�����j�jA��!��3߼�m�"�MNl����H(
�Xz��$'�Q1����[Z�DH�u!�!��(~��kI��uB%���Q�T�c T?|�(I���^]�+&�!� ] j���4O�mNYk�Y����"�8�XV%'%�Ex�7`	�z�)��u!*�]�(�`h�r=Gq��򚎋!� Y@��iIğ�F�Sd���pa`^O��������+�Ŀ烁�6i������fs�	!�K[]}���DpP��2�ܐ�=܇^<#*c7�����b:k9���a��G�]�LU��6�'�?� :���e�$�0ӂƔ����� �9T�r��=7��5�CCܓ0�7�j��w�z���x~�P#@�H�V+χa6幂��;����=�ǈ.��Y��̕�қ;�7���̒sA�*��`Hr�:b�}F�;���]���߿1������9���_.@�4�"���H�D�FҘ	iŃ�L;w�ה�t$ժj����;@������'TXp��ga�M�[C��]�`AV�/O�PF	�ir)Q}������䠝��x��N&RW`�|}���vEk��������WϯIN�b�Z��������s���k��7Ve`���b�#rsBƷ�J���G����I�l�I�3��b~e�� �bqv���¿=C^v���,
*?���qt+�m�z�UHvh���I������s��K�K92�����RB���PmhK��$�JIz��4�.��Y��w(��y���4
�6ޝ�b�M��
�|�FdB�K����^p3��E( P@��!����FԱŃ�ց�)1"�{m�F$�|�MDׯ�x�_�>{ �ئ�h����N젪��%�=���K�n�$X��
DSU9Iz�f�bB��)6`s�%�亍/�&�a�ڟ$m�Y�2ס����,��WC>��xmp��D�eD�%����{Y<��
��gb������keh�W�/�����T�c�(Ѻ�l�.G�lȿ3�cն}���V�Z�l�J��e¼}�~��W�[s��9�L�2����K�9�n��pu�m=Gp/$S2S	Z38Br��
����o� WZ�k��~�$����X�n1Z�l�汞��5���Y&|�SJ�D�F�*�H�P@"��Q��X��xy�}��HXΕ�J�x������B��J�a�~zbU��Ss�`h���⨾	�:���k�fͲn����&��`��k=X����2�T���S`��E�	FO�K���4V�����P3kt�>H*c������d7b�����r��GI�[:�::���+�
�b)ĈoZK>ĉTex{��26]Ġ$L�.��}��䚸�.�]a��P��ր�RJ�����(�J�n4���<D�>}�![���D��ߙ}�3������o�$������Bi����W=RZ���?�\��?Dlf+4�8a�h�mΏǐErә��ȡV݊L��?K'W�e@J�����8Dt[E0W�#�1����t��î�BR�-��{����)y�E�����G���f��=�E���#,�U���m��a��.)l�GOHm;3�}R�V�'�U�2��y�A���s����bi�q|�5~��!��>: �17]F�/��U�%v�'�o�-�tR\����(̿&���1x�i����s���(��G&r!��l���7�F�E�(��!�ZGu
9������iGg���5?���i��D�]�.l+�Z��ƴ{z<D��1�d"Ľ��|M��`�2���gYŨ�M�v�nbu��%chb�wtl7�l���1ãe����6��/F����L�i�Tm�GZ��s���\�h3���f�k�K�~�2ǆ����P���S���|��}�_��dy��N�;��th�9��%hu����^�{�Ə;���5�$`&��@2��C@a�'�5��%2�q]1��q w������`��2ZS��0�����%9M���70��)!d:n<��5�ܣS�o2^�	���/�8xG�ak��Ȯ����ۀwM��ZH�}�ǆ+w-[1���پ�-E�Yʂ�-�?�t`}=~�,�����!�5�R|�@�j�w�$@����H��,q�Ǐz� ����b�'�r&8��3(���|����P��Po�m���V.g��W������^�j��N;]w�ux��>�8h��q&ʸ�͚�k�p��H�!r�cwx��$���WPS*�D��)��?f�I�����FQ��)v�蚲t;^O�|�&�ݠ%�2,_���P!K1M���/��g\�/l�:���W 1J��j���$ĻI��C��	B�k#�ՙO%ꟂV�t]��B
M��,�\K@�|�҂ r0l�!�H�aQ���<���k�Ou� �h�����x1��7��(O����L���-Ξ1�qB釅�����Q���ٯ�49�5{��2)~��-u]�!��O��BC s��k��*����?.�Ɇ"@"���\D��گ���"�ԭ��N�~�Lr�ot����l�'��KlZ���i�H�T����~W���fW��"m]�FK�lt�]�]�)�C�_���#��&�7�o�i����>�O(I��Zn��A�K�Td�\��%��]#&�|�`k��j��¤K]���a;�ơ��P�:ҟuY>0�"��3�H�u��d���ζ��3�x���L���MV�Ē�29nb=wv?_k�#ē�>���E��ue5���е}H�a�*���LD�gw1�/������0[�b;�~��oW�,�(}�f>����~H�t2���I��U;���#Z�g�O�ۻ/1O�՝:f�'�Q�9�� ��:��&�����^�z��X���H���
���Uʢ����:�9X�a"8\�����r/e"bV�A���T2LMt��:c{���i1�Ef`�Z�b�u����-��CK���gh��>b��*���V��np(�`y�q  ɽ����=���ȷ�m�M;<��� T;Q'H�h�����Bup�BC�0+hA�������� t�����}�/�Q9W���Չ�Amt�vbD?<3�9��+���&��pp-!�(��ц]^��<�ˠ6r,�p�qH @��I�C,6�;�a.A�~������̴�B*�R�b��Ԙ>���3Q�\�O^���E��2��nU���<w��T�qU1�D�Hxy�_�ȇ��2�'�6�P�ʶn~�����!I餝JnI�\�6X���R%��੻��|_@4����k�C,𲔬ִ���ݲ&02����F���J�]B��(���sr
چ�<�w=s�$��3$�+�=dz�!E�G�dm�/C�f��x�����	MGKPE����+z&�u���?Y;ܶV����(���LL����\/���5��s���m�I��#�7�����iy4�+��\�A<�@P��T|�ܲk�Kk�wzVXo5S��w�g��uY_i8�5�y�f���ҠQ!ٗ�}G��pgE�^��TE�b����qG�ƹ�;�yHp�b���;�1�h=�BQ��T.�x�*��I��5uez�g��p���b?~oe�GO
(����>���FD�g&~��S}
-�23U�{C�~X�ל]����il@*���A]i�?�!8B�(�Bc�0Ͽ����e�̪�!lS@�����O���M����]��;��& ����|�1mU��C����{k�����K��;;X�ث
�îQ\#Z�c�������7v�>�
��M�JV[E�C�s�����z|���[#!Lߕ,�f�t��n�\������ E��ZS�vj�Jzv�m�Y0�.�����=@�p����+�3��?qJ��n���
��C��i�]��Wӄc�J��q�s�hy��^���fsЃf���$�IN��V~���Rs���/�9R��g��iA:r14�q%_�7�k������+֓5s���JM�?���\ u��B�~h����'��k.\�Υ����f�ܘ ����9�%������N�ҕ���)��.���9�q�}��1�
�2v
5�ĥP�/5� ęVRA'�Fl�W���J��>#�c#y�� �q����>"��������|��0f��8/͉��r�w4])K��t?�c!H i�c5�>��Š8w�<�%[=�ۆ�@a]��((�;U���������#Gb���Do��
�Sߡ�zY ��t+�i[���$ʘ^�S�&��fB�LV�+��F�C����3�+q����T�.� �����N�4�r���2�~Ԩ7���G[�zu�����0�뺭�p�z@R;A�'�r,KQri���ዕ�/���7� ����'gw��ޚ]�
J6�eF�%@�,�o�����3�g!��������k���1'
�����1R�΅&���� ~�!�	�I���P�'�%���2���wJ*Sk�[ÿ{!��7��4v+j�h#$�xq���� �`Ƙn��9��N�m���:�Molk�.�_�˼�'��C�dzt��Sŵc�/�E���	[���|���j\zF%�����>y��tpK"�uW�4��DAt���-p��!��r)�]�|��:͆��\%�Lޖ:��w���W�0A�}Ul��!���|��&$,3�{�%�����ۃ/%�'Z�bM���30tV��ܛ����X��9���S�|Sr�n�6H���E�,�Eu]����
|�E��3�=l ��)� �Y���xMɢ̚rSy�ע3
��-�����)Sp��
b�F�8��"߶<���u�[OB9��λ�"}g�u���<6�ܸ8(=@��Ԥ���!!��.����2i�Wl�+���Z��wi�t"�S�a��("�{C�{�*f��hKUh�kW5�����ܦ	W5v�������@��¦Q�@s�x��6���̹��i�6Fz ��)��XG���f `�?l���[��D=�ˊ��PZ�5��aq&^�"�������f��ߖ@s'9�&z{
�bt#Czz�	E��pnsRu;_v?���(��������A|,�^���'y�c/B�K��dr<xC�8۴dD����6[Ԍw�ͫ���ׇ{c���]a����Pꃡm��}��%�DZePs6�ZǗ�\�X?��0�9Y�'1��;������^r@X�S�@���2�㴦f��jB�e荣ڮ���ǭ�8�-�� �MP|����a_>I����F�K�<qCTTy�����V1�qA��%y=P�#[ P���__o��Y:p��.�]�'o��j����ԗѹ��KDm(�b\�ôI
֬�P"3�6 ����v��V�5ZZ���u�f�n�lD�[|����>�e!���̌��i�0]mC�2?��j�$}�K`�|Kk��#B�(��~�?$^���ә�_�8X�d��W,9b�]����� �)�Yw�p���krڅ�@~A��G:'aGp��1'6�wi�^�2v�|v��GV��P�~�#7�-۾��w;5?-������eaKS��z���!�KW��%t)�#��V;`�Yt�RQ��(�k�\��e���r}�$�fY��W��T��������O���	�au�꣣s�Y���4l�9�T�A[A��F�:�;���ߝ}�m�q��t��C����/�_NA��޷�Q�l۱סJL�� �c�����vTʳ��\�#X�V嬙h�J&���S���q-�D�~�8=-1#+�s|8�~h�kW���xL��m��z��>���6@ڻ�VL��D^f���9M�h�DTc1K��Z��n��|gpZ������D����A�NU���J�c�_`?��b
������(_���x��cCq�7�q�%����^��ݛw+1��XI��?y�R����Oo~�j�Gb�S�(xF��zg����C�4��;�pP����v�uҏ�(O�G��iu�����©kמrDf�O�NU����&9�Z��:���Rd�3U(N��Ⱥ�)���c�e��m��O��H���u�T��=�CH�{�����ht��8��tOK����pJ�R�z'�VPGȀ������:�.�۞�f��Z��_]�Nm@���6���k>�@�A�4*�<�Y$��nu���"s>W|@��O����E}ZǦ�q��.0Y4`Y�*�B�I8CѰl!�vH��e
�1M�9N'5C�=XRl`�?i:7�8+aC\��M�:�8�
�U]��5mZ˂����IǺ�.?b����=i�p��i	���w[�S��y�����9�20��cN�B�!�%J8�����ob� /��s�!6�d���J���\��l���H���$@��\��}ݐY@"2sT��fB��`����2�祗ߊ���2�;F���� _IIHD:�B��')�/�*�Fӳ6AvRQ2?��]������&��"����F�Qz��Z�5�%��qP%��?ú�_m���H�]�Z'd�������������P� ��|1����m�:a�Vl�}���a��7H�Μ����o`u�D���kz�P�4Q���Jx?
�+Ê�/L&�b�c�*Qr�<ǎ�"�i���?9m;d+�&�|��������B��^��~�0'��2�/�'�����٭מTJu[La���u�7 #�����ǬX{Ӄ	�1�p�0@���ty�������Ʊj�����l�q�Ԧ���S*��fw��I%�߄ĄE�x������%�Μ��?I�X�&�>c&к��X[��0�_�Y������+W�ĴB1�
��e���˒��'�j��w�6��·�0Ɓb~m�xPg_la��L��"�P�q�Z����kL�~UD���f����ou�]A)ҡ�Y����D���,!�}�YJĥ�mh���/��Ŧa��ד�Zz����E��f&e���7кoܳ�����ߓ��}�R��i�}��T%m=|0w%M��5+���A�C�b�'f�x���!9��/|Xk��!D0����xo�q$�Q�U���(�{��Pu���>�lRB�d��*6��y{a� �1�<�\��_��;�JR��3�O�-�7�:O� �'�nd�7�������޾��u�n<���FKo�
v�$���=� П�:;��2+�U|�˧�v������!�P`~�>�4���6���n2�(�5Y)�Q���Ϸ.C��*)w�7a=.>����ȫ���i?�u�����&y���W����j�p��$c����f�'}�"�8-�����V�e��ۯwC%��1<�y�^9̯A6i�{ܮ��k�nyd��o=3Oe��Un�#�y��p,�}9BЌ`��Ҁ��Õ}���;Պ��HA�����	p{7��E$�s��%�Ke��ܵL[4�s�7�(pyY]6�ŌʽU3�j�{���^d9H�r��s������?�,0���@�r�c�G70���B[ϼ�i��D�C�Tx�n��&@�99i�D��2�6ઃ�Xy���;Q���7��)��J!��_t��`M(�KwN�;��2}�����f����Jb���M�[@���',g�#̠%��'A @�� ���r!t����_��q�֓`���,�C��^�;�sCs!ڊM�E��kg��4Ȭ�y���6q�<���U7��Ly(�����' ~�RjUbe�Q�o�2U��&��P�����^ Q��� 5���j3D*�*U�1�:��{�x��r�%���#M��A�v�*�K����C e���ޒ�B��߂��ac.��h�װ��Ƨ�/��5|�b/��8�h&�2G��L���N���0d1�܇)�-�z�y	ܙ�L<Dv?�q��>��W�a,q%d�?�J��އ�]C��Y{�%��O4p5��<h�=�&�ł��M4�q��9ɿi�h�h2sE=�8Ġ���&�ϭ���&����*��̘��Zo���6c�������oC@�tJuu�n$Ǥ��������z��2F����x�Y��f!Yu��T����i�U�J���4��$_����ꄵ%�%� [w������C����+]m�6h!o���.B���C��v��;����J��8���cGF,��Y_����A���f��X�2+�Z��W�ӈ��+�sg��UP��8�6����,�_�(L_��8u�[�}������?&�=t_�l�7B ����DK_G�*�z���S���
���	Q����d�	��ٍ��S"K��I3)�GƦ\Ր��0�Q8��5â\�*�h FwU��GTD��Q��1ʌ��jiͯL� D���[�q�/�kᷪ��gM�
o0�I�O>&�Ay���g�;s�}�b-vAf��,�F��N�{���&� �X���P�sܼ"Td J#���JG�wE���빲�u��X��b�ªv�]��&L��$]�k��j���s|�	i�Z���MK�=R�8��E���Iͥk�2�2�P���H��i��d;���#u��&�zL����u��I����bEi3����p6]�`��bFul]���ȣ��)h�HAfix�l>���)���	�Ѷ���F���X��ǔ��`����JtA,��J,�� _��g���r���?��a�ԎM�QѦ��%9p0�R��֟.0[ĭ��f �6I@i����#�C�c�kJDIx
�]�=%%��p1EZ�P��vB��q�j�j��pP�&�V'2��1q���:�����U����4r����[�6:������, ��PK�c���o�~Н�VX@�W� ��ʶ�7B1
����6&�Ǥd��I�n]9e�R~H���'��\��C�f,2�*<�J��Ykj-Q��"7�B֍�X�B^d���I���(���&��ٌ�e�͙��Do4WV�����Tg�A�jR�1縗A�	��8ea��	s���	�J�����H�g�0Ӎ-q�Aߕ��8��s�������C/rő�������t91C�D��c��|�Hʘ��ǋ7�~���	T�0�l��>�������e�Hn�*4��:/����9hބY�i�I�*N��]є<���$��`�{�O�U��4�|�:��Le��J��y��mi�7�ZYHR�㰿y���~�aiR���3��t� ���V����a��s���g�0�YA(J,��;Ͼjv�J�	�y�#�:��0��	O�����*��WuK��K�t+J~��E3FaZ��	n����Z���c4�����/E]Ȥ��%z�?ޞH�5MtC*��4�trqO{�ڻ�fqC�?8���#h͈����EΚ�Ez:�.����Q��"���ܒl�c��2-0��('���rt!�� �M��q�k�t`�q�B�]�a�5E]�Nt�=�B�)g8!�� ��?���1�B(J����Sܘ+H�Oe�)�Uu��2G�xb�HO�-�Xہ��`y\Ayv2���u�"L��qC����ݣ"�d/vY�5�>k0RiKY���L$�X��=0��� ��٤M[��˺E; ;��h釸�Cx�iX0; wF�2�����|�)!>�:bd~pI�C��hG9�X�f�8]\�T��:��0@��g�
'�xiJ��ed�"b^>t�u�Q���g+�d"sE�R�e�o�%�,���I�že%���[�xTW#�MP�m8��D�tTh��lE����Mϻ]���gm`t����J(M�r�Q��zT�̍G�
��k�cg����sv���>}�E�䁫���
�j�x����^�,�jNU�%����З�V1�	_[6t���~��������
���c��At�Lg��,���̮�N�wD��Ԏ�/����*��SRsC��{��I�hw2~и�''�2�iV�'� �p4Q�"Bo+�T}\!��s �%ah_�xS�dvP{`���+�E�e�"
���5$t�GP�q�o=;%
R�a�������0�g��'3��G�de���4ɠ,��&�"��` VN���OP/�:SӨz,���/=f����ˣ� o�*&D�gG"�)ҕ�k3V����y��4�"�˄��aD�ZV�q�:o2ML2�'�2�혂bTT��9�W�\0�e���ÏA��Q�c�2v��ۉ����JS��&��&�-3����x��b�ljY�9�� �[v����jA����4���5"{������E|UY�A. ����]"��[:�����=,S'A�s�+��Bu�/�2�$�z҂4���.���4�8Q�������{�h�
"� O5��3���]4���\ӫ�ƙ�T����/	�Rˬ���	J0+�z��Rt�Zɿ�:�I��@�E2o�a�G�K�߸�i�9O��#�d���^���[ۖjܟk1-�S���Ţ���K@�Y+�^p:�²�6�5|׍2HEi�)�6��<�����N�)��M#.B8�=�8�?PP�8:Ւ�gJ$v�*��*:� ﶀ�t���{FL;�p^>JW���t�P:�Cݽ6\��*c��^��0|��L�������X�nj�y{%WC\�f�(;3҂�@G�D�N���>��>���s��Z��Gl{�';!���Nc�6Wǝ�,�QVM�^�ӝ�69�V�텶��H���3����w�O��ĢueXj�i��g1x7��U
.��h$ٲ����6�EfL4�����+&n߽�~�������2c�:�8e)B-~�I����t���K����Y+��UE�w6v�E%g��<���D�Rqʆ�W��\�3҄�hon��Z@KH�>Atu�?�<ۿ�;����Az���c�}B�X����l|NV�cr�)>�4z3q.n!���u˱���m6�%hT�m�����ƙ�)k�(���]1�t3ծ�.��(J���Dۤk��I)z/,,�ro$�7H���V�(뒎�t���IĎH��).~���+ ���$��&���!�A� f��l��-u�.��0��G2�񃪪'�C��4��f�=0p̤zug-��s�+���2m(��ֿU12ÄS�i(�c�e!FN٦�=ܥ���aC�}���f��]�AWҁd����P&�f�۩�Z���m��%n�灷��Z]���o@(��vB,|f-��>>��C���_N��e��{�^�,�� 0-��^�<�r9���]h/"� ��?�����7���K#����5�~��c������N[ǟ�O)��#�Yz�!�����w^
����jݿ�F&vLĵ*�ɼ�UK��o�%�\��M*�h�V@����V6@����>C�C*���{�v3�[V��1�b�\&�t��U��JMhq�:^�'�t�uH\)�^h�0a	�{䑦�ʨ�"�4ᑗ_�#22p"�.f�a!�N|�e��	wtH��cͩ���vw-b��A�M�}���6��W@Q`b�ں;�&��ʀ���p�	�D�UW1�3�[V��r�fbq'��� dUa��w*�'0�,W��*ͬ:�q[��!�PDj�?��|��,r��g����O�<mp���D,z5�!k�6n�!��S1�1��]���=de���u��w]@��{-�v�j9ۊ8�[8�c��8���K�⴦�P��t� �uBWS�͌U8)]^���'"�!��mS�ϷA8��_��v*��`�U�,"d���1��FDȸ����L
�I�����wfd�7ĚƾEK.-���*5��>�FFҸW)�Yj(f�ˆBH���Cy���K��^Dw���L.��pDsNi%��H)��\�X��L9i�
�4L&E�lr�A�3���э#�.����Yz��IJ�]�F�1)i��5`O��d��ŷFV��� ��~	��R��"����7�_}��Ƕ������!��.?ǩ�S���v��ZÅC���v@q)��^���9�*b���x�+����q��"�����5��m�䗿!9�{�+�疭s~�~v|�Z��Z��s:��i&	+��<��S/�%�,��(�i*f�?W��/�r���h�9��2#
!X�8L����-�,]�6��KfB2M�EGJ��)���������:�]7�/�ht��a��x��R�A��u˨�^��#8?���"Kz���Qɵs��d����
6hg��-�j�{wuj?*�c	!�E^U��D�-/_�I��DyY }�}&�O=���mbq��>��!r�����E�xح{���lj�y��"#�|E���k�|�=S�Ϸ*�j��:;d��f�0�N�S���7E�lRz�&������k��z�p%m�0]��8NОp2�W��8Sr,rw��� =�Cj�Ű�<h��M������O8D+=v�T1��s9�\c.��J�p$+��F�etX�X�����}a.���������2�f]�0[sU4���ʠ>l����&�]��Ng���_%���~��A�{~��M��з�Hi��:hW{Fo�8���%�.2;��i@<Oh`I2���J����X_�/��@D| *aF�o�69O��\�1��mp�A�V���5d��������߳k�N��B-�>���}�~d�R�\��%4#�!��/W�F��nJ����|5Y^�f�z�'�*U���_5Ǣ�:��?�.�_����1��;k>@�Lr���>��}ˠ/t�`+A͹c��Չ�y�K�ǡ�brdx�t|���ӓIN[��X�9�J��r��4��"�/P>6�� �oH����ښ�;t{R7�7͎6�1�L����۾$��e����R�t�c�b̻=����'��`@�*4��b?�.���BOt�@����@D()8a^U�aa����Z-U��_("۾��1�Pl�D�T�IL%�e�Z��(�L�d��>�ڑ����^W�	oΨ��MP�i�t���@1��ִS\D�nn��#��~��^R�8��/4m�"��+p�C���<����j>�o�#˱_��{�����%�H������:�{+w;[u����X�H��x�sv�ɜ�Xup�J 'm����$�y
(�](��u��	�ay�[u��)�k�f<pE%�r}*A���A|2�҃�6�S�FH�؜ǓeL�\�KWw#�F<SZ�
�>�j�
j��3��C���f,�Qp����B"���Z�IzP��`������Y֛)�#N=e��z�P-\���Ɨ����'h�߯�
�(d�Lk^��q+��f
/�N�P�����׭L���.��NH4	sc�Γ���na��G�/@ZR��vJ��ew4��(0pNZ�%%7�o�������6�^�L' Ck ��/cK�Ñ�`-���$�\Rx�� q��0\M.̌Q�����Q����o��C��p�� ����� �}��(b���]���)D��H�o���.���꬜��'c�~ayu}�h���R����l9݋�]E�s��(�)i��mj��1���rD�a۪��]�0�(�
fK@��&unT�"�-cïH��N�~ ��1~�6)خ���/���iN��6�M<y�ll�7|wr����ڸk��퓯�_���B8Ӝ��gH�
��i~��+F\�A�l4k���2L˗�c��Y�Nkci�*�"����pp&82�} �#��ry+��:"<[P�A���#�bG�;/6�х�	<��㱻��Xkh����p?�/J:G}����r�["{�ϫ:�T�ދ��Ԫ�7���{��HR:˽3�$L�v�&
h�!��b]B���Բ\L�/v��Z
�lsG/����K���ѣ�K�2Q�>����A�I�[.ڌ�1�ˏ���5M�d��C�[�jl�98^�i�:�}%Tx������p��!#p
�q����s��9�u���X{R�4
XG�����z ��2a��^� ���+�|4�����m�˲�ͱz�s1�.�7��/[w�è��[,j?#���Ig��ϟ�)��I�z)�Z���k��t�ಀ+A��X�n��GгF��P���tp�#n)���n+X�=�׌	��Y�:�:����	҈�ТbU4j߭1�7�������R��%ȑ�:�8���-}�R��_��C�B�)o��J�ec$�hdA@�zI~�@{����,Yp o�8p��C�ev��L ����yU��l��N���%���;B����Й��;���N�VB�[��ɓQFM�;�ta�kH�����:��*-��~���;4�u�/`aR��cb�ՖB@l����މf�@�t�@��s ���/���&ڬ& �L̰�R�B��%��A��3�NIԡ{ڎ.^���S%Ώ�1�l�1JU�,�������P��*���
-tRH�~��Kb�� �aM��D�8>�-Tz>�Od �g��AEf�m�=���S�O��䑀�C��|&o��7��R]��D�C�	^�U��7[��s�G2�����Z[��Kq��ɀ9� ��})�"�r�۸i=���B�����mE��w����{�o�k
�XԒ9z���m��!�W�T�#6X��iJp�P𜧕+���g����wt���Mc�DDw�'pW����OaAE�U~ut�F5��[�k�"�������K� ��¦5��_�A\�A����5�9�p��|�N�Pku_�����������bm�_^������;v%nm@��.kh��U zp��{ݘ+&��!W�c =�rHŖ{
��B��� ��54�#�
j�� %\��1&�y��(����Y�����I6�oZ�.��p��f��SE]�@�Խ�u潊꒔��)�IQ!�m]�(p��zD�6k�	���h �����v�=��t��%������Rڦ�zU�5(홏U$&"|r����̄F���g Q���@��-t��w�4I����J� k��s�蟏�ɀe����X���{x�o;��W�f7�YP��tE_%�J�JWb]�,\�KO�$HCno��r��C���C
76�)�N�bJj���yF�����^���N\�/|ə�y��%��]�A^Fߘ��&5#Ǡ�ҙ�'������rP�3����QH�&�	�)g�nlf�"�}��$m_^l�)�#��s��"�*�jFɓ�i�=Ț���8���QJo׿���ػd}_>����D����9}[R���l_޷Qk:�߂)�~#�t��8��C���Cƻ)h�m��������O��r��a>�����16yd���/�r��R[��(�*�8t%Y��S�r�FR��=���a[��P��)0m
�sT<�(Ø�,V�Ϲ�>rk}�P���@Y��x��04���v� NX�!�nt�_�Y5ԙ�.XS�u8w���p���a	�י�2�6oڷG �h�*
��w��J�5���9����T� ǃ��8�G{$�q����� *LRO�X���z����Z8�$&Ϫrz��XW�"�,W
c����B��y�'nj�?=ե�;�	e��ZKp|�����Z��'��m���m�@`����2l���_=k�N�xĭ��:ݚj�B���ԑ��]���fTp����9I��^(MF]G`v�Wk�W{2:�3��Yd7���qvM���0f;Ǌ!�(jϜO�:>_٢���Y�L�ZseE��3���!�0�;���7p��_��x'��q_Q� r?��9����+�z돒m#�Ks������G!�������-��[ᑴJ��1�OlqHW��)XO -�R	�)oo( �	;��)>�`�0��``Ѣ���$D��F�K�Q��NA.��*^����hQѼ ���:E�.�70sXRT��YqYHa���n��Q�n�-,�W�g�;��u%��jo�S����&���n8�:#��q�E�i,@N���S�T�N1�2oԥ�<1���� |�^��E�8g,l���`��JkM<r�Ƿ��a_ŅBɞ0Qy#�}"�=�d	9K|�/�:��>�iH�WP��fZ1��`z~��WY �!�VQ,��>	�{��+c��EG�?bI�a�CD9��?Y��Lӡ�:�I~�)�3��,�X\J�$LA�u:����?����ń��Q1i�4�#.*;
8�@W�]�S}�b뒿����Ӟ�@
��Yn,�o�" �4��"���J�㵫���5=���?�T�Vl�#�}���1]�m�H/C�v�ַ�����b��Lb�c�e��.�K=�Ҍ������^���<h��U�3�J��kY�
U�L���f�ۢ�tįH�<ܐv�[n^�g�HB�N��sA9ؾr|������㩏¿�2����p�?�V� �R�A=�įL����ۊ���ݻ �)��{̄��EV#�h��`1ykj����/sO�-������j���	0]��Nx��]Bюږs�P���Ξ�\,P�y;��)`l3k�r	�v����$��Co~��I%��c�RK�ۯt�C�j��J�%i2����kW�^s+��Bq�G�$jD��!x�Չ,�C�Ĝ�$���F-6!��l��h�L8��OX�{gbo�.,�SE��#�Eu.��p���)�\�ʗ�Fگ�%v��/G`o!�ń���aKn�Szsר�G������
`�)Ƥ�]���BIGi�܅l��N�g8����/"ŻI�HUP��_��'Ji�Eu1�`���b#yx�/���F�s|De���n\p�'�@��Ӥ������Op�af�f��rJ��g�l%F�{���L_w���-�WQ��ۏ/�M�S�Ҁ,���=�n��IO�|�5&�쨄�q��@J5��-�"�B�F�9�nS�<��6�X�&O-�+¢ڊ2^�<\����������s܂OS6~�����CJ�,gXIѳ���SN��/c��@�9�S�6�?�E�ȅy�Ή�Tp_�d�-.>�����!J@���,eaT�b���RI���)�񩵅�����S`�%�$�_��mkhC���6��8��(��+�L�i�H.�"���^L�".8UAmd�����x��<+K96�oY:uU-�����`�r���*��2x��n[)�gA&�׌�d��[ &6��d��M8�?�'���q�N�[�W��V�`f���H�jWU�4e��J��n1�Ed��E@pӣ1p\c�Ě'`Yb�WB͎/=�3��
��}��I�s{���5���u_67�0�
6�w�֙1B{�����J^GPK]�E�U�i�;�FE>@�[U#�,$  8dJ�1�7��Nfm�+��A�TJ��.+w���ic����Z�wH�;��i��x�{��//� ����!;ֹ#u`�0;D*�٭�Z1AR�m�¦�4{�F�(� W_�X~+`xV�e��d�W�Dr�H�-1��HR����y�o��<��y��t���z�Ũ�Ƶ0|,��
�=M1���݊sd��mV->�����T�!�9�'��2
9qH���U�����+�E �>#�!6�' :to7��4xVê8�;����/1�ֹk�<��t�"2���aB��F'a2Q:>��Ȅ��kѝ��S��Q��A�'bT��8� ���m��>��� 5Gc1Vm���u��e'���:j���F�[�d�U�X:�N2����b�vy]�{�HE�(E�`�	�q�ZBd������1����R�1���6�mbjP�)f/܃�����PKH�<Iϧ�
��D�b�t+�E	�H�Fl�M]�#�ZvX'����gn�u(�&Q�ͬ:�]�Ƶ��57J��#�Vsl8�+��Qe1�:�o/��{@��0�g�R�}�����Y���y���^]��3)�Y&8`W��7��y5p��k�"���$�Ҫ��I�������I��[�I�b���������]�nNtK����U�I��������s��N�bJ�
Į�.��ō?/���^ız�|�SR-ω��Rz+p���mx
ֺ�Mjleųd//�v;ؤ5ᡔ��������
1�_��u)���w�����e��{�M�T��5��gJ���˵���=?��TFч��@ �J�Y��+yV���<��t�0��7o��`~]���� 3j��B/���/�bw/� ��(����#M��k::�
ݰ0H&�:m�غZjm~��~�s���Ξ������Z}�5��dOq��Hhl�I������޹]�"�삇��g�_}C�V_���$8%����-�^���aD��x ��Nm��4FM����Ta�~gi �Z���7^6�>�܏��|?M��K�!���c�3�z'Bڽ�R��3�^2W�<b+N��{������W�P�X�SES��'Y�0��1ԘSR��Lt`���� n¾���8?6Tc�'Y��ZڛzkI��3~[
��!'���V�K��z�u�=H�+W��D�@����y��GS�O. �V���Z��!�����w��+�r@
Lu��Ȭ����Kѳ�Ĩ����7V�/W�	Wj���@O�v��LĀ�d_� �Gj�2�ėM��3��ev�l�6�����8�^85#�YD�;���P�

s����l�:N�?��
ú�(&F2l��z��=r:,s%-�4H'n�T�I�:�>5f@�g�F�C�f���_�HƩV�$����=y�'/O��tt������U��(.� I��'�U� ��pl�a����q"f7����O�f^
EE+qq�#^<F%�&���r�T�'^U@�n�����׽G��H�^mM��#�l
����8�)&!���3ġ[��p��M|2	q���zf�"���pŗl�_�Y��a��_� 2����SI��]�U��/�y��P�0`��nŗ�-Ø�u��&��^��^F'�s�3�)�3/����_��iϵM��,�97��l�
�7���b,Ң�ig�0D���I.VБr8�&,�M�P�$���Z��3�I���:2C�fd�\0,���)wf3r��M�0����}F�ǣ��^94��r���T��?���+o/ ���+\����8����E�	�J�	�W����W�� �^i?=��! q��0  �>�O~�����ɭ��!�X��5J������	 ���!w�h���Dϧ�k��d��V�_!č��o�(���&.�6�𲐻��V'UI�@��՘Щ~�5�c�GՃ��]���TNh)�}���Z�>�`E7l�X���M��7���qs�䈕;���]��5��<d�HC���ƃ�F$���y��y��7z�F}��Ec��,g(
���RX7lE�}�CuY���= �o�G�������L�*UA�-ζ��)�+Yi�	&9�A�lqN�����[jE���K$��HzJ�F�Iʷ��ed�-y����������9A&�'��_SNVƭ8q�d��=�Ӻ�N�:�*	CNU0=9��9��ފt�DAd���:�
�^��g���L��0�l�>��lJ����D�4��ٔ��?�U���Y� �����Jjuy�,�7Y��)��R��^S���F�=r� 4���]���u��L6�kb�Dʁ��4M��{A��p|������K��]AE�[��1���r�	5��SI� Up_�s5�2�k�6�1�Z?��=��P�)�W�1"5e�])i.*�ITڹ��E&wp��؛�,�$��D���e?^�&]� �r���2�Fk�J	��L��~�h�����n��ۺ7�`x�/0	y��hq���;�jױ�9tX�B)ݗC���9��*�s�����J��Qv9	I�u޸�-1٦�M�w"�"��]p�~�Iݺ�c���q����oO��:5� �&-.��PNm�l�UWp�O��xUg�U@������@�-�oܓb8��6k��E�M6���O�B�[������I�?m�=_��Z5�0� �����$��\p���R���m�b���P��8�����%wA�,�ziU��5;�r	 0�O��xM�{�D�bzZ��\{@��а:�ְzs!��=���G��霥����Ib��,@V��zi�����'��W&Fs�"�<:��q��B�͘X?�)8�>v��'5[��}��|���ꮏ8"sַ������u��-�#��ZX�F�0�Q5��@�r��>�,J
C�6&��p�%�$�����Q�����(x3������M������܄��B��m�Ŧ�"�E�݄H\�?�j����zR
?Z�SL�w�:��Į�4�+��b>����}��3l�8*�������_@Ej��=�b�k��|V��S����s�pl���vw�C/��/ ��-��,*3%z�ii.��4F��׎�!����pژ\�JR��)].[��I%���z�MciWvu`����}�J��w;Y�6��Q���BٓU`��pUߦd̦���'��Ň�Z�.�|����a������11a�Q��¶+S�&_k^m��>�q��{�Up՞yA��%0��6NJ�LS3��eBJ0l��Gy��t��E�CT�
q��bs��e ��uW&����"���0�W)?2�`��cː�a��5�]g6�:C,���}w�6.;/��K��%��҆����f��kO�&x��+ �<y�L
�;xޯZ_�<�mMLq�p3�hW��Kk�Z5��mł�V+a-иv*����8SH�ʈu�9���>�_3J���o�{#n-^\\��ߢ�A��
F�����Ks\p�0C6i�4��I���/1�B։��>�@Mv�ȎL�٢�-M��z�߮�`W	V�� ٘l[�l����q��k]2��k���N���:ܝ�_3�k!�Q3B�&��NiG^�Fnţ�R�N�j`1��������&�:����K��gjL�m�GQ�4�خ�-�	�y���,��_3�o��&�t�E�<r+*%�!�&V������n>x�#=�t^������A��e$������O�0�K���[���=>��ma��:��.���z��X��(�E�˜��=�1�^[�IG�Ҩ���L
��؊�gg�6<�D}�=�3��`ߪ����i���4�C��8�\I���_��%Ym��jU6� '�̌m��Q�g��o�Y�f�hO����|�X��5�ّb[��ޣ�����`��7{,*����q(S��uS�C����C%��.l��������}��P>��M���,X�Ƹ�r)zTq?�����h�Ŵ�F�;g�v��_Ku;պ�_���"ʠ祴��,[���0k�[���S�0��	�(���5E�=�\n���Zk�QD��������FpVZ�:\�Q�^.߃ꆧ�H��g�n�u�]�^*]��3�ͅ����S�
�.C�����f@���!7��[�H�.�$�$l����[����S��ptrQ��	����nb���/W^�:��f{(�?6L�)�f��s����	��W:/0��ԥ���
P�T�װub�@�l����18y��	�޹`k���U�V�F���Kku_��G�5;޽�	�}1��-P����w�^�#DU<���$���}#j4�]A�<˃�@��^��O���?jkv���!�*Y��:�=*����'�2j�Y���8g�#6�Cr�y��]�����2Z�I����)�=�3��
�9�W�v��l��		��|�|݅Dە��U_�����\R ��ES����EÊg��'��#�&�V���*]�\}c���:��!�$���j�5�F�xt�Z�5�D��d3B���[ii�3���0��ҥuP�&��p��oq���m�@�䒢����O���z�	�OK�E] E���-���]��ҙ�ײ�Q��:uZ)��[��'U�:ĎJe2������A<��=j3w��4ƅ?ՈDzή�\"�ڔ�~��	�Fs�N�z�?�ݠ���,��yF:�}ɭ�����vp�������0��p��&n4���!|��^ˁBN큧d��D<6����uES��D��Zt.��9�,	���DT!�ھ�PD��z����Z�[c����(o���X����ɡ`�QQG�)]"p�����4����a*ܵ"�e��FmU��Y�I��C�ͭ��@��q��6�Vx׶�R	r�[\��ڄ��b����@f5��ҽt�[��:�m	 jsu��Y���3��쐈��B�v�w�4�@��Z��nM��m0���g��\d�1ώr��u�w�������桉LW�����*�8Z)�`d�?����M��a����70]��F+�4��K�����6�"Pg���@z�Aa�������Sz�:�,;��Oa3RF+�/i�E�:�|�0^��/�D��h�#mÎ�>���������R�ɦ a�g�~����6��꼎y���:�c֊uG����v7����
�ݖW9%��[���M�Ds3ld+Uc��=�a�^�"��z���^���h�ZM��>��<�����-��s����S����0�{Fx�z	[h�S���ɦ|�s1WV$x;�����㴢�����������h��@�����2����5R OK3���e��Fr��Z�:�	
e �G?8hd��29
��?�V�W�2��_���[�B|[�8�������9�	R=�����j:-�\�폺O΋ph�SJ'����+���|��O�����M%��g�A���8��^XK|����]Jr��h�q�%o�'J����J��4Kw"��L��z������w�З]�u�.3�G����Am�j�Gw���7����!�Yl0r,M�2A=z�>����4!j�'����`�`G��VoV�!���C_�X�l���2mV�Lw��!ѯ���君X���)���PꚇrcpS����-�w	��e��ԉ�)��˽1��p�7j��Uz:�=l"d6\�2�ⓤq��;�Ŀs)mw�*��pD���^*���
.��	a�ğm}�)���B�:��)6�e��(�|?�r�h�BUj�:�(����q�mͧRs�<}��Y� p"��?O^�� K�%�1b���E�c2�jvI�����Ŋ���G%_A�a�/�9�e����II�A$(��ͯ��F,yQcᄅ^r�@GDp�H��hC*v������$ �_x�&��1R�l7/H�wZ.m���Gh�c&��;�=�ƈ��0��9jǡ��ccn�Є2� Z�O�#9�	�S��������>�7#ȝԹ*��In�:����K6��~�.3D�g� =]?�����#���4��]������������m1&�치���:"�?��o�k�Jp�V�_��QbD:��ή'��:"c�z�sϴ�y�B��L�&B�j�\,a���|r	;[�$���7ϛS>�9�/�g$��  WTH��.s"�
��Y�+ ��:8��ɞ��&С���e1!�32Pe��F��LBϙB���K���v���1
�-V�ϖ�IZ���L�k�:m���Syj�&;�~uA��a�V�y��,���B|���ȝ�&'�i���4�k���.��O�e^�:)	et��¼��S�N��Z��6�U^K�Q({�_D�c���2���a����)y��|"�j�����LJB�$�1R���x�8Sx\5qo�I�x�5m�%�e;�����Y���\�ܬ�jS*��>&���o�6�h�K=��N���,�!�+\J���R[`�W����ba.��w-,���g�d[]|����S]>�-�Dy=�8 Y�0��:y���g���.�8؎dEJ��]6~5#�&#ӵ�2��������>��(��!}���7�٠��-����q)?�7����`�@�X������ Y9�K�?���}]S�)�hD�F	�o�����8�/�cC�\����ZaU����/���c�ݩw�����G���x\j�D}ـ� �k��+4)��C�rr�.�����@���um"���Ow���
�]�1���SF�5�S�edX�~�(VZ��&�o��5%�7M?���(uD��M�W4�^�.�R�=^��~�r�)��w'��	 �z,1�Su��xveo�F�Oɔt�+�
^�S
�m>���30r�tK�-,T�MzT���ȓ�βNVA:�i����y��x�ޅ:xN���:pM{��Za36�`�t�A된�>��9	�yI�]�y@��%�D̗!����f]�*|�1.�b��1(,��"=�,����/����|;�qI��B��i;hx��b��c+���f/ps$���G�z���<+�+��O�UG=��4���A;&�y����ҹy�	�f鼓�C<��g0����ޱ�Ro9���������$�o����|�����#����zM�VlE^�H>�����rN:3���<��|�K(��7x>�'����k����G?�4����:k��Ck��,RD���O�L��QJ茏U�e��r�xF|��6(e�:�U���o�z�8�]�6ǳv���'*��?�ѐ";���K.�"�
~o�x��۟��^�45;8��Ex��=!��]�s�*3�������`�r�b�\��sr(�U��1܃�I��n�;O��IOx�������:~�ju�`��X:Xg�d�w�/��>bԘF�1F����jx��X��o��kǀ� ��&#DȠ��K����2+*�ڛ�3�y�,��x`P0;U��;��.��E�s����q�ӂ��eup�ٙl}J�چQ�MQ-����c[ۃE�;
{�x��B�
�Sd���B�C�����)�����;���j�.\��ǯkc�p���r�-�Aꚨ�)��"�H�#`*��/�=�L.}v�2�9��!�Nr�)�ya͠����KR��gə��[kV@��8"J^�Bo�/��(����L��ܪ������ye�{�X�`�����9�ۅ�;�G��7�k�Ҷ
���ps��g���&�.Vk�FO��S�{g�..�1�hd��%Ť�SBx:�75��b[yK���`+z�A�R�y�Z�	� ^?���`�}�[�,��~�̚,XT5�+\���\�)
�C>
����6-<X�rZ��f��X���~�w��T!�5����X��Q/�Pp�=Q^QӦ���/W�&�ώ1I jp�
�7EW\�e�s����<�('S ���O��,��m�G/�n1v<}=�?׻X��VP������Y �;����������0i���D�I�̨��ݨ��;9���������v|�R�#M'Iڕrc�9�I�A�d�p ��fbȉ�#CC����2���肢e�Vt�=�R&�C �C#�d�j���aW�'�f����[y���IE�{��W��Ť�+����P�\V�8�� #�
��!1U_�~F$�Z�;7�Mv��eUcaF7R���_�}`F�c6��x~��ϐج.��9��(]�H�`�6��ҏ�^,�t�}
j>���f��]S[�� `��]�K
��8v��CÍ�����y�}*��,�t�E���~���o��I.�\6G�����X����(Po��A�ז��T�"~�]�x�&�'��t�S;�Ye�,���n�x�����
_\������C),�B~�&�]�8�擯g�)���M��2�QR�[O��76�	 ��d�H)���D���L�|��&Ƣ�L���>(V�q�iu���;;=d_ݣ�
����C)mb�k�Z��+�m�:�]���^v*\hв�TC��E%��T��A��Ex�W�7s�U�Mi[��3�N�����ŌKz�hL�]΃�X�@�G�\ĉht�߂�P�!&���H����X�J�)>!^qy�¨oSO	�/v�0"3ju�x]���s����; �� d�c����.�!�Y��,5��� z�ârΆ&�v�s!
H�Ge)�|��<���<e�����>5�
A��cVΩ�0q�7�Ss���X�m�Z�@n$C;}B54������r�,WK��Op���"����I��w'o+��9B<h��s���a'�;��d�aӗ��D4�n�76��qk�E�n{:���t_i"�ϴHq��=�Vp.�9��q>��6%�����"��*�W�,�?1~i��Q��\i������0�����̠�Q������>H��Y��ܺu�� 5(�#Lk�ۈ��ô��bm�wC �����bE:{���T+�w�1�Ä�`�� aמ0Z�
b,96S$�����I���0���k�`�7��͸��_������h</��-�P���2..�r �����˱��'0�J�w���4��Q�����H@�o+Hӭͅ���d�{ٟ]�U������Q
f��֬����&�p"������{w�^)�D�<�:��uL�i��� �~�QQlX���7H��6�4M�@f�\"���-��w���')�����4����v�r{Ƃ����eE�'�K"�]����'5�l�)s�M\eiB�n��9��Ly�wG���k����)J�K6E:�I�+��͏��$I�;=m�5fSp�s^|ʒ[qq��NĞ�_?�9��l@��pV~3l��Wc}���?$ħZ(��Kw�%ȕ�9�ަ�\�{����0���Ӄ��>O&b<.��DԚ����jʏvP*��]�Ȟx�� �?n��v��{d���2ލ*��+������)�n�d! ��S��Ya�-U�#�|�UY":tz�+�<oCJk�b��V�Se"��D�<
����y���e�ˠ��g؍��o
C=H�'�e*�L�Z�`��+��'�-,a�H��g��OSyq��U�O�3nTc�o~�M�H+Щ!tN��x��pj���Wg&�<�?�x)�poD���A;*8�g ٦k�������s9�3#Xɿ̶��1(�O'E;�y��ϒ��,a;�p��V!��vDrE�2�ah9ن����~��.��+�%���4��s�(��ݛ�+*�y�A��)v�/@���>AW�⯞�0:%��;��0��h�7�<��L��?29jKϛ����c�UӞ��m�=��{f%�i����zD�|<�M�2��h� �=�����u�e��LX����W�:@t�t��RG�^)�'��ߪ����v�W/��.��M���}�dC�]��ߛ�cxE.��_�Ҏq�(�,���<���3����LX�g?�}�4`����	���O}�����Z�B�jR�O�:�
$�9�c^���\�wi�I0�.m]95�92���pP� �Z���;q}��|��Kt�����)��'ܕ�^(�Vx���+�k,�y�M��U��p�d�Q�RxϠI�_��OP1�S�?J�/��'��C߅Lt��0����&g�P��P�*\���gW���X���`�Xr���Ul�s<~���`���{����e�I�ő�d�ul�iD��8�J�C�t��NM�T1�e�}�] ����,�b��U3s��2JdZ�x�LE&l*h'|@Q�}���F����g�,�*_��/� tK�e�-MH�Vw!��"M�_Lk��I��p�L&�>�4x�}����*�1۽����˶����1α�� �PN��H9?K���$�f��5��ep�#�Y#@���e�=IJe�Yr
�;z�G �2��|uL�Ꝃ
��O�9I�{]�!���F8yA9��
V!/�Y:��`�)V��f��k�6� �����?Qun%�i��*-L��~��S�SDg���"��X�y������C<���F;�-K��!�xh��
��EpF~�bыVP��!< 3؋�]>�^�����Cݽk���XFr5��*,=)�D��t3q��v��<l?�����' ��}�;��������Qo�`�hB�Q��0O(�s%%�nτ��/I|�ߤ��]�uw+ЫCy����ч������|� V���������Ⱥ&���g���㠻+� Ã"(<��2�^�3�m�Q�"O�ָt�:�zj��h���O���[�j��Ia�`V�/�T=`X#�WP,��n{>/��:I��v2�����=�D��݇	u4�|�!i�m����L2��U��8�Q�N��I��QXK�?>"ծQ�*�4+�=�����lYN#�8
ٗ&�de��+����:�ᘱ���F R<��z�n��zhZK�p�p�.��	!�+���zH�U�� 5�3,�F}��jdy�j
`���zfΰF��ԛJ+��d��y/	[��W�����J�M!̩'
�u�E;^Zl������b*S\�kIn>��������(��fq�aQ���S�_,�~�L����K�I��`�	']3��@�/Z�FN�WrR\,�Q}RR��7��?��2�c����`ˉ���f���t�.���2�MRvM�
nfj�R��S{��fX�

-�Fr���P�gp�ﲠ�i��gn���;ISd�8�^���4K�Щ��J���l�mٷ~6i����6�k�*��\���r�!�[B�������=�~w��7z>�o+�/23!��A���W�2�L�9�T6:|'{�ڮ��^Lz�z$��e�?tL��*�+�)��Do$W�d�;�O#d]��^�˨ �Ic�{%_x� ����![� �^=�b��E-0G����,�����<�e����W����j�.�IT�o�b��6�0���C��:&{�3a�C|�σ��Z�t��i��l�vC�ų��&i�_����C�ĥ���ᔐ(�*I[��WB�̿z��%�����`�"�s\��M�R=Sf�c�:<��ĝ|�SU@�A��6*gZi� ����<q��=F�D9��ծQ+�*�f�δ&j	���Z'��x\P��P�� +���d�34�p�4��vT����	7W�b"E�%��.�Q^�6Iب��2�%z�Y"+c�$�*��oj��U��P� ��i고R��n[����4����N��h�-����*�8��d��p�*]LM|+wl� �U?M\���qՆ܁����+�)�k��(���J�̗��׋=:��
�!>�Q͉vB�o`߷����baZX#;M�J�(�v�,���~�K��YH�����j֠�J ��\yo�,��)��<���]P�r����y]��:Ҝ����!�
o�Qf"�C�X���b���x�P	�1@2�#
�}V�U.�~5�}�(�UC���0,^������-�zx/�Q��|	�L���̳��; �a�k�>G��˰�Tm�'�+��:1�'�I���,�m�������Ѿ"N�Ε�|Ԅ/�+
��*=���:����#bi�W�ِ��.��Y����Z�d2�4��9%:*��hWUo�/��5��1�}ᡤ�,��-) ���ݱ�T��a��܉��x��|�e�<9xLM]dv�g��مI@
���I0(@������A��lX�ͨw�W~x�jh���6��(�b����1{�q���jIe��0Z��uf�N��,Xi�Sf�Ȟ�k�	��3z6���?��ߢ������shf�m	<ɕJ�]�&;Uc�-����r`�z4�\�j��#\�!A=���� ?�z�����'��F���!R!��B23��&�� Y,0�t�~ت�iZ�gh�)�@��e�6���)�a�j/F�^���:�F�U�<���	���T1)����R���o����_M��h&d�V�t�1�depXlT"`�KW)T�jeEg`���J�⢍[�s�R�$|w;�D�y!���l�ؼ�KN��D����~��#֩
ċBw��y'P�&�,��(�����?�0Va��Kp�����TOD��Q�K-tͼ��~O�����7�7���͆/��f|�`�e)�̮�9�A�W�;-i�;�!s������G�M�U|�/t�����=ὔN��znh&ԳD�����Q���#L6GYi�����n�� �:<�U��o�n��S4�������r1��q�ނ����w�<U�0]b���,	��%}�M��OS��Q�ĵ
X\�J]+'��Kˇ��a��$/S�����p��ۨ}~5?�/�D1�N�ja�7�
,G.�{�0����]1�gW'�(���z|.g�;�/ �:M1��G��:f<�����M������ڙ�R��7��	L%�آ)i��HTN���
~�;c`��HW���!?\��g�����'�{����樛�U���1ݚXT�� c���1�����2:�����\	���uZ�
y�� �$�A�ڈߔ����#m�e�Fl������K!_��%�(��Z���jAo|��s$̗V1��`��p������������YA��H���"�zBU�����#��
�U '��DI�8@:̨�yT��]|����|�|f$N�i�ŪXd����zd���YczZ�R{՗qܬKD�Xac�Ho����f�s��_9�f�2�T�B����
zT���VK���B�|T��U�ôP�^����1.qyRT"g\�J������l��,a�;i%�-���:��K���� pc�A5-�E%s�x�����s�Kl~�@����+�evM2Q�PC��!��0c�����#n�<�FR�7���}����tE�-'����_�)�Ϝ��ؓ�I�OL���x\Jz���1������Z|2���8�zY�_E����O�A���v�Ϋ�n���j��RަS�9}����dg_��y[�On�ѧ�"E�Gs�.H ��yY�0�`��-�|	[t���ޅ1�6��/�{�1)p��Y�vq}l*꣤��7�E���R�E�ش䖕b�c��N�ޏ��5IF��˳ K=n���A�Fg=����L�L��� 6�ev!dj_g	��%�R��p���$$3Ƃ?4ށ"){l]��b�@�!5~�G���xm�q��Dl�aWR�ҁ�e^��1�0��
��YV���4O`���[�A�������&1�� �<MƔR(2X�2�FJ�)Il��Uha�X@<���8�\�By6�·�)�LX��P�D	�vϔ1e(��<g4��-=��0M2/�3 �(�^�ǮyA�2o��^�	�&m9��[��ZŊ���Y�*�f�:�Ҵ����|��BA���9�����T/x���l=Ǚ�l$�Ҍ��y���t~b�� ���k1Q�f2_�IRI��?][��0�Z%L.u��կâ9O�<��T]̒�|�B���?��&���r���w�q��<�/Ȩu8ʤ$W�D�R/����[��EBN*8%>�`��|	�Wx�Ӣ���'��q7.����bq,o�R���eoJ<]�g�����2��Xs(V'b� a��yՉ�!�Q
�B��3�YTD�ܺ����2�Z��6خ]�tQ�eG���؅|?��`��e�+�>a�JQ��]��7�IJwT�\9��U#8&�n4N�Ny��p�@�!��X�W8���al����+��m�mJ6�x�gй��|�$�4�R�[ �l����l����>w�s�~�&)�I.f8���3��ø�ɶS��@/�Z�)���Jh�&��T�V4���Q��d���%��	��9'�ؓ��V��,+�(*�u�������>^��aPB�[m���٨:�9zn�����m<�O�z���G!5�~��{"�OL>38/W�v]�3`#��ne��S�d����CE����1�w����{2k�<���`��|~&�q���p�����Y�\<Y/~Vxv2_}����c'3�ķݕʖ��[<��7ߨ��D�OW�!H�^[��^�3��;�8�l+�Z� 7��������
X�Q���j���$�n��̝<�ϲ	lX7�gm�R��L���'O��U�t,�l���z$l䍼՘��`��z��vc�r!����@��9*J��z4�$?Ƈ�*`����w~�q�]���Zi�Dw�r&�/f'ΓL��ZoY�}�% �d�a�<ɲ�z�W�oi�^��]�{�zw��4$��z��j|)��=fM�B�Re�H�֜�MFv���w��I�$M�ޘ��R2�;�*�1�e;V�ܚ�֟̋�,�?3�7in/r�L�ʱ�Re�\rZ�/�e&�daJ����A�QU^�854�$�J�9��Yev�T��aY����_Q��b^�CB��|\k'�A!������\mp������l�/V"o2�	g��m��S�����pޱ�o[`��	���ժWx�
�C-J׊��Uv�~XjR��w�����y�Y}��.��#�A��CM]�%z�5K�����Rr������!f}�TO4���0Cp��͌6ۊu+���^��������Jr�S3٫�n��+𔄣��il_�D,wN#Nu�bT��!dr�=�������q��u��+���<ֶ��d�V����#�������{F'Ϙ׫�E�?���S*8M�S�N��M�(D��]�J��<�I��;�/�	5]�*�u-� *�v�Ń�v�=�"CȒ��6�'��'!��O)��U
Ú�7�3Eo�C���/i���NH�����a��Ē��B�Kq� �Ч�J�b�]���O�è����D�6Hs�����n�8��Aז���ᔓ���P_M,٩G�%�x@e-���#`�)�U�15K�o'���|(�B�b�Q5T��΍Id��'d%���{�[�˶Dɞ���3����4�q���ŜS�0lV5�gdE̐��u�03���>�r.�ў'��i��0
���匷�-�h
��L*�6R�d��*����N,�HC_����y���h};0sȹ���_(PD"Ύ,fA���嫓�2֝�O+����������Y����3B2��˪��wݑ`���(P<�G��_����[����fo8B�gN���/�G�VU�9%�Nu�&u�#l����N�@B�!D��{�q=��ޡIeM�}�����LB�G~����8����AJbJj��S�f%Z�hK�а�
��o��v-���@��?p_�x����z1�}ٟ��g
d{��@��6�W��"��� +-�I�6��p|�b���^��=(�#4���L5��hOiBkw}@�_��VFQ��� �l�k�`�B�Hɚt�h�=���+a}��ک�ow�%��j� �q��nk?:�%ۨQw�@��;`���Ʋs9�z7&e�2��x(�~3r|�m2�寇�1��GB�;�5����=� B��@<�Q�__k �3t_�����[b�QI������7+z���1�¿2�!���wG���? ź��Z+��]O�OW��cfJ�������e���B�qyU�EYJ��q�;h�q������+*�[ (���
�� ໐+��Ԯ�����5PO5�D}����IED�h�9��}��ҭ�Y�e��fA�iVL��W$�(�<�t,�����|x" ������7��he3R��(�ޭ�KZ�9'ZE�����CsC��Z���fܼȊ��l'�<�䌀�̛G�e��޼o��!,�sKX�M���k\�&p�)�!!Eh��/FN������"�;SqE:R:�xY9o��l�%<� �x�C.�ޢ7��� �}�|x��|����oOq�S¬ C����)9Kñ�қb�7`�p����aN2L�/�2��J������vt\�M��&��M� B�u��%�djD!0sW`���D�.7�}YVI$8E8>��lm��w'���CM���?�g�u�l�m.�9����+Z֛���h$���{��]����^_YǫtAm3p���f�Z�C��0�E��"�6��"��5_��ML�VF�HuqI�KIYz�x�G鿀��u`���ٰ�
ȉÀ�#���]����(�P���Gg�Wc�wIr��;���Q"��T����ȑ�5T�~��+�����v��k�� M.dz�h?��Ϗ .����H��Na�x� �ü��4v�J��^fMV���d��D�s��ek���� Z��%�;�N�9�ϊ"]`ƹ��Չ}���g���SX��ᵥ�E��-�Hc/�J��N���J{PZ.�5�cƮ7=*x>���I�IͧBj���c*�Fő���.�����ٸ�ؿ�w���ڌV�"'�,>vU{�~�T��9J�p�L�V�|o�^)�!PI���o���C��Jo_��1{I��@�>g�R�Ll�X��+���%u�k�>�|/�~����Ӡd���D~�|
��£�$ik�sQ��+|�%v�VL����h��F��q�4����6.ʝ���@������A��/wW"�J8hƖ�����h_��7���\�;}�ձ����BĨ�.�?�ۯ1ò6o�����M�+��"u��+36;m���L�Ň ������_��p�)��e��޻��o�l����Ȥ���SQl3�	r:�
5V�ޯ?f�A��P+Vbn�@�pAb��:�.�|�O/Ӡsi{�v�J��Gŏ<e4A�o8��]�1G���#�}��+"|�5c�B�A��qr��K��u���(��R9�V�5���G�#cL�3,�z0���G9ޚ;}+$�Ե�H�0wOѪ�#���UC��y\��m�3����fYoT�K�I?1]�6~�"��+�mf�ܦs6�$�5�>��ȋ���C�5RӺ.��i??����VO�a!ϧ�~U a�Ue�傽sӘ����C��	cڏ!7�1��h��?p\�w9���\c�񥻼�T���TQ�*u�w).I�5�ɟ��f���:!��t�Y�rϝ �w�{=-o�5H���v���U��J����*�GV?�������/	�c�����N0�U١�h��L�#G�����B�?p�}r��>0�1��1�HU�:,I~�C��L��
��2D0��P��՜;��Z���󤵪��PZ�����6,}��e	I�³�(,�6��x_u��A��Ҫ�����(���~��z��;<m}���D�B�z9��h<,M�7�J�߄T�.��d�4���ђ��m�L��7�1�S�� �m��d�< =�$�5Y@��,9���܂�H.�V ����!0��i�i!|O)v���M�_y�)��K�V����-�WB#I�b��*����-���̒[�dH�q�b��e7�6z�?[h ,=�%	�b�+�h�D^��l!��F�U�6π.��~��q������
���Įd>����H��c0^$4=���Nm�~  �n3��6�zK��$:��6�L-E�}�W���i���!h�J.HW��U3���ă�t�7=9'���ïai��*>�qQ�������y�_�A�t�{�1�	�o0�l!����
;�<����ׅ�&i�/ߝ2�z�>
Ȝ7$A�o\�I��(>��$�1��z��~^���8� \ˉ��}N�ۢ h��0}�
xH%�4��9�������#��ݿ�P�d��>�[�v̫�
��m�c��.C�}|Tu5�@��՛k�(��X��oy.S~ H�iv4�nC}��$JY��S����x;�St�1B�mCэGi8�׷����*��˔sQ;���YYڬW����/"t� ����\bs��+�)ƹE_�2kx��Ĳ�Mts0v�_�!$�b/��qP��K�Ǳ@���8�&���+8��@����yވJF�(�.�[�E�^
g�9��?��q8���z�lg�m�$�M��+��X��b🛻�en70�����sc7�l��e�nV�Ҡ� ���3�Z���m�?�VQ���X�2���pO$�ThR+��Ǫ�Υ��hː��7��Nw갣 �%59��1�k5�ڦSK�76�wb������%�a��{_e�7hm��Om�h/Vm�l�L�T?xI�����\n85 �'�G��eo��"FH}bx �`:���]�Rqn��ƣR�Z����54�H&��?����I{Oz3�&�`�m�D5���sG{R_' ���	댫���C��_��7�[�\��(�?�3��64q ��%�D�Z��G˿�ߊ�d�#&4��z؎ԉ���7�n6½T��+�y��$[�I/��?F[aSt'��n�*��ea�i�	��w���L�D��h��KT6����s�O!�H��BH�k���{	�r(>8,k��_9��%�V��Ƚ���f)ԓPl�F���� ��� �Sb��~��J�1N3��6�"� ���9��R�
������~�8�m�\
�1�d��h:H�	s�[��[��J��-��Pz��w���<6P�fس�͖+���5*	Y���|E���� �^�;�LO��@W��i���I #�̸�7>8�+���>Ӎx֢�C��\�ߜ�i�/!�1��X	�4�A�>I�d���#���$�6{
�ɳ�Л3��:��pTD�]&$���9؉��.0a� ��� �\��Z�J����{J3�����ÿ"̤A֗6�+�G|ǜ���IG�V)�HŃ�7�({�#˩;G��)��
;2�c�|ll�򺫔�-ҹGMs�a�Q�[������& ��bZȰqyyt,%�R� �Y�+� �xOT�ʽ�{�i70����=0�//:�0f��(&�>) kK�8��t\��N6 2#=��j�T.L*-K ���avD����~=�(ظ�|ߎ�N3i�8խ�
����r��)��S�E�,�G6��iLW�"{�*�G���o-C`i=)�s˗�MI���{	.�'j���FBv͵�A�oj+�7�R=rPgB~������u�QS��Ô��FRcܹH^�����"�[�������VI`�=k���
Ѻ�P�^.�=�Fѫ~���B��<p/����b�D�jV_z�F�;�����)���#C�!����7N^��2)v�xEGJ� ��[+.�枨�k� ���
�L�}�28�q�f��r5�fn��gn���:<���,c��C���w����C��&z����óv{�Lr��#݊�8P�P��|n&�L�!�z=cд�n;�¨dVr���xgAh���N\1�]:m"Z\��2kћc��?�^������U�Z���8�Q�]�G�M]@n�ʺ:�r�%�%�f�M�J6��=�� ��X���\2���d�8��vG|^7�O�q�.��_A�ݯJ�l�Ζ�4������#m�f���h��7n�\�^���,��,S�Rq8z��攢��]�{�� ����r\�F�i*>�n�����{a��hX���d�zt��8����Y�3��Ut4�fp��T�^��{߳v>�u'm����5�:-����?�\%�x���"� �����3<]�e�4Dn=�v�Q��
���1%:��i�p�#��`[,�$7}��LS��ь�l�6��4N���r��Y�֒��%��L�{�s=�I��v�\��*�rRb? ~ژ��ߎW��z֬�*�M��(�"�:�[�7��2�ן딗�9�#�����Z
�s"�R�]�>���Q��^�xy���F�f�i������� �AsP�*7�v~�64��M3kӚA%���i���'�CK�:3����~/����J�7�i#a��8�������:��,��w��J��+��j%�;��H��f.�C�Twǉ��L����JL�e�X��b��BE2��#o�e;1��·x��Wг�@<X�%����I	�4� %��{�#�_�1~ҁ����;/NE��/���m� �ِtt+��*���㽙1٤�b$I��z�%�SY�� d��uy+#K^�v�V�7m#K�\�κ�g�̝�G08���p?ˆ�_&���E����:n�7�)j��_`�z�}Q���gM�����޻%T����-xx�7A�<�;G9WR�i���F��+��ڎ� �S����ļ���n�ҧP�O�9��``�s^\r&{-Th���EN�u���AeZ�͛sg�)�M7�5���z��gy����y��S�S�	���`@ם�ka=����'2@V�9;{����e���V������ۗj�v[ ����Q�"借�R��z%`�z�K�L�Ⲗ��h�!���.o�H��U1&�"סF�;i:U� y_mU��k���t�v�h=����[hC�T�{.�ɞ^�5H��5O�F���va%����R8f�KR�ׯ��\l���^��t�.J��o�!	>qy^��%�{q�-=EWڏPj�4P��?w°Mf��{��g�L\L�b��y�R>J��?�$�5>iG>�̔2�nS���������\q�Y�Ĕ�ٺ2L��QE�(!��S3�	U�$T�Y^����I���>0b���oyǉ�I�������c@�!3�0o�pgx���8�y�b���я:x��U�PEN9�I���;gv{���^��3wqYv��P
�h#D*�]��Q�b��E��Ʒ�����;����['�m���(Z��Y�J��s�+�����z7�(ѤL��h�R������̈́�{Ѣ�ܮx/�w7)
2i�}�ܣ�����QW�CZ����V��3�-<�gY@�C��.Qe���^��5���o�*Ȯp�Z+X�衏#b���+�9kN��r��_w���3������	��}t�zZ%�{%f@�!9�{?&ġ-���:��*�"N��8�l$^¹H���Z%�?��UӇovXhFI��pR����6�+<Uή���w�rjK�vQg���ғ�r���&lO���ԑ��9�\���u.�ϐ�L5�;z�1m1N��|�4��%y���j T�c	ۘ�֥%��,ٕ���� �f���~sk�P�Ow+�V5����������w2���Nm�X�����\�1~���Ή������X��V~ϊ��4T��S��)��.$N��E�~�SB��ۧ�y�zbG�6��g|
�Se®:�ߢ��_�k;N�K� ɂ���ߣᬘ�Ѷ��EA���C@�����k=��7Kez����IZ Tˆ5Y����#�g�Y�-_!o��$I�)���@Ƌ���߫�3u��1 c�z��Va�o���iV��tlF�y	�ه���8,-�g�
�T��R���۟��0jo�����&7 1��q
2q�/,�p*xd~�hɚ*U�ԓ9� �mѥ�T8z}�������z��=:du4'��m����ܝ��x/3�,����r�p�Y���͗b|qfeN���	�2�&K�YC�Q�w{�l��pktk���:T����gOz�E��V�������P2�Xs���c�a�r{&�ɞK�T����
V1D�\�gMK̎����`�>e�w`
1����-��E6��G�)K�Սq�fX�ڍH-d�Ա��w=&�"�~�M�e�;X���vt���SFb@P����&�4�T���'��/Y��:��S�|�$���%Z��"�jS#�'8?������`�vC�;4~�'Qc�ɵ�q�
�l,:�`3�
����C�9��P�YϷ�ߕ}s���s@����w��V���*��L|U���+��;��N_W�\��F�i$r�L��F�ͯ�ߕh��43�Ӑj�JӜ�;��*J;*6߻����a��?�>�c��g��ds	6NUm�;`a��::���(�<�FW :k��n��{��<��,Z�AlN����_�F�q�����:Z���P|sָґ��$�P�
ׁC��:�d�/f�  ��o�{� 8z�
ezʺ�!�P���Ť��5��U��P��B�#���+s]:�)�lSg���Xx>�-=��(D��2^�߂�pH�7�j��*0�u�X�����;F�F�A��
j�q�XZTgu�쎱eDh�ٱ+Ͼ�q���́�?�����W��OG�w�T�Qg���6 I�n�^��6�A%��������e���4�u��!G)�X�@z�i6�1���g�_�&��AM�;�����*��fN��a�W�P@�<j���6ȇ{a8\��Io􍒀���^Z�7;�˄�:��+ԅ�����sm��D�+�Gɹ��z�qk�ODH��l���O.�&#���j�[T�j�D�h�M�	�zo	���H����W�8�E�.O�&�"�CJ��ɥ��cwR��&!H���Jn�#�Ӧ�������8z�j^�~�.��N�B
ԩ���k�9��J���h�cL����	rr�^c]�F��~��0���Vm0`/6@*?��2U r��*<�4u{��������/-N!�~���0�}��m�߯��igm���&��K��2y��>�ބ��q�4~��ஈv9(w�8�n	DD����@�D�T�7t6�OK(�>�z	�?C��۷�r25X�؄�;�|��O���%��;=��ͧ#l���<���M������	*�A�>ꐴ�?
�M������{_L���m����I'���ܻ��ZŬ��6ԍS6�q�8í��(�r?$���� i���悯��vZ�%�K �n=Ǝ(�4Ѽ�/'���k�~`z����lu�^�yDZIBb���!�cͮ����gA-�m���R�h�dY�p�] �H���,��7e{o��Iͮh�`&�Z����9#xܱ�e��)���aXR3�������d�sȜ]a1��2/2D&"N��8�T������T*e��^w��K@>dkT���� ?��ca��*)\Xi�B��/%o���{��<mK�u�TՀ��v�Oמ��'��(#0來c P�E� 5�e�p��Ӻ�c����)��}�<~���_<���ol}?�[�[����)�Iuo������=���B�:��;� ��0d�}�	��0�����<�H��~��j��d�4��_�6G�A��r�Aecm���p��ϵ�u�:��Qj~��gٰ�5.����*�?"k�){G�'�ʏU^�[RJ����K{���4'�kH��Ωp�l�i����|��B�nsQW�(x�V������:�]��G���!�OO�����Fn<��?��E�u��/�	%����@�1k<q�d��>�pn�4{�b��X�P�g�OF!��|]j�c�(�OX)?<�f��#2�G�O��	c������+���sŻ����6���͠�+Jj��S.*���qw=J+YӾ�b��YFF�5�V����Il��Dj�0X�OkWߪ���||�X3ĩ��L�J�Q�c���vS{Bf�qJi�q-�0�f���Ve�$�	9Jb]�+kW��ĝ�&�1aC�8����b�w�u[i��3e���%�̤�R)���� ��y��[���8ߩsE�0,�W9�b��v��W���M	���N>2�<�߮G�ڹ�XAz����r*תt���Q@�������r���� �i�HƜ���E�ĥ��*�ƨ�ؾ��t䳛�[Zbx��DR�V�M���&�+�F������xV����
�&��"C�iw�(�~���w�2T������w����$���ӛ�Q)tni/Ȅ�D�Seb�`�m7��oC�D�(=eI��p0Pݚ���h��Yk�zx?G�פ\[��}ߥ����_������g´���϶Y5��N8���(Rr�Vd�k�7���4�� ��C���|[�D-���$x��:�a��=���������Ɒx��y��v���.Iw�������Fz�r�X�6�g��N_Yv��ŴY��=;��lgc�2���B"�Gu��ͯ��R����mG��mYC�fUPs�>
J6��E��.��-�~ j/�xYqY�G� ������B�K)12�a��c�=6��p�b�;H�3�U!�$����'�U	b�dy# \R��	$�/3K[i�;Mﵖ hŖ]�LQY:�aF�񆻔n/B���VêB0ҿ���8�a	z��D#3�9���Fq]��.���O�4�b|�wr�ۣ�}�ҹd���I�Ĩ����^�_k��Ѐ㉆�`�.�4�l��ys��$�-��wp-|�� 6Z���v�0X��rd�C���ݡ��F-��Tvۋۈ��|�%�|��yn�+�i ����#Kh��A������]"	�����"��B�	��ad��a�_e\*^�dVZ��	5��E��l}B���9E�U�֭�L���o�΢�A-w�~2��J���7� ����.>d����F��m�k�ȿ��_\L[�1�}#y\�<�G�Y-�(��6qMp`�����_�9)_�����/�QF��ސ�W���ѽ[��R���LlZ�DD�,����-c���'���?ax�E/��
c����^k��B�SW����%����.��~����uS��KU�~�����p�������h��O�>4��)�Ѣp�]�����4V�D6Vt%�Dg�V��� ��ϧ�ߒ�ҾK����XUg;���L��QpC��$�R.�� OO��@Ԧ�+k�����hP��
�5?M*�*G]w�S$5�\_N�т���i���/�f��>���x����u���~V�x�ɷ?����x��K��QՉ\8������RT�.�BW���4	#X�iS吗�\��=�����R������샞r.Û8�a<�.;�7�?Q������(u�bZp�_?nu5�p4���¯7����d�����Mv�aU���jX�p��ױ���"仪|PU������[�`�Q�f ��% %�8rFS����ɾ��>P(��C8k���]�A�a�c��J3�gQ���,�	�������|�$/�0��vHĜJh�u䯼IC���������E'V���eͦ0a��[=R��r���!y]���:LT�׸Y���ď:�!f�:� ԨsA�<�.�8rT���$3�����"��� ��K�~�� ��M(4�q.��#&�������g�gӣ�Ú�[�H`T�d* ��$�SQ\0�2��]�U����hgNY�b�D��R�fʇWYx����8~�e��9��]�{��Dph���u�X�:���A�'M�280�߰2XS59%I��Q���;]��bc�M����
HS@�),%bw��a ������g��'ʇ�
 	@iV��Q�@���i��S���jb@�x,fDt�&z�ԱVW��Ћ�����Ûtv�V��S|-�4�y��P ���a����~Cހ�ff$b)H@!#\P��Z���#��|׽J}>�B��k�Z���L���p�}I�S3�
5�Km�$���O�#'����k�e�[)1��^��k���A��΁`C�)u�SM@��j���2��m-肃�̧j����a�9�aQ_��5��x랒@.6�B��ǆ�x�..���KY��P��t�$�!������]��\U']wq9��GN8��v�Bo�nQ�։�k����\���B)��;��
��{��6Ĉ�"�Xn�B�Ԑ�+�I_%��(V.��W���-h��t.#���gL֝�+���*�����"(�V�@��E�=X�x��
��ʿ�He�W�2���R&(�����Bҥ���1�s�u�	�d�ơ�d��3�A@J��D���?@U���E���N�w�I��\��j���!�����Ã@_�;lM΍�����B���^7��W�����ffÉ%ԫ���%�Sx�y��{+���וfC����!T8�fsw3hHl�-����MTz�_d�,a[>�i�Hvaa�ۄ���=�w�r�xé��V���ͲYE��q騩�~�<3��q���%~`� �P1¤�wK�FzQ�p��Zá0��WZ�iPe���/#:K#N�I��۲d�<��8`��*(xH3ױ�9���T<h�!q��eB�-i��;�8�0�Ny �{�C�Z�ع?�.h��R��Q���D��t�n�#�tH��N�`ḹ�I����7���DIaJ����XF/���~��@5�=�j�}�yE�w�u<��q����3P�ˤFR�a�׀F���j���Y�j�e���k���;!}�O9�~��󲚣--���Q�P���F��:�DfL	ɪ��bʓE��z'x7�6P��''���'��!��?��훂U�1}��Z{����ǆ���2�'�?PC6�� �=�+%�������;��5�b�΃��R��u�3�N>�ǘ��c�߂�6�U+��/���	@_��jm��h��G�v����q�?+H����S_ɫ�>A�
6��nx�\�$p$�1�|TWc�[�yf������vx����' �L+�V�Ĝ����DO{n����x��8��N~��gtOБrX��㘣��@Kjw'���yR�G��n� ��e��D�;B��?}(���ϛyO���w���5Ⱥ�~���	v|q��`]C{Q�V7z���iVp��:06��L�Ն7'�H�3�h��迨�#��ѭ���0RX}�|[ئ�m�Jl�VmC^y�iv��pP;��z�5GP�
���Z���/y��x��i�#����Q24�X�A��{�%a��ǅ�{�����h�����~4�_֝P�$�&�0G1�휥�Ҭ5�Ы�M$�:/�K~�}���(U-J.{��ihu�2iA��	�	��2Hƾ˛G�^��af�۱���=�o��D=<5Uh��w�L{Vؓٽ*NE^s�Z��w0�{�����C_<�c2�m���A;r��y5WC�0�[=��x���;�����M+����v�bM@6da���=�Jѐ���
�\�����|A����F�$�����3�=�\K�Y#��8�p�e"�)��r���
 �.`)��f���*�S�0db|��7�J��.���/x#��L#�%%���+�	��r^�i�]��?�Y�O.�L�.~/�e��9��|C�G7^��<�"Z�:/z�OPXv�I>~����٘K���3�x$%"�6�1׉ӋԫeѨ,e�X�^F�X;�ѷӣP�Q�:�MH����%�'Fr�Pd�V5ڊ�6)�)<�G��$;�@>�m�!	��0��+~MPD��
��r�m@r����Xٸ� 1�B+����зЀNĝ���\@��+]���:����j���X�$p����3�y��8V�c�Ej��^���D����Q�s��Z�@@6p�Tz����5< ��)"��x
	r@���k�=���N���Α�>]��`�%}��Ǩ	���{T|Ifw���8�%�İ�c-B� �Z�Ok��2�<�
p��E91y7m;��T:1�e p�gF�Vϸ:\�Z.�_�]��Z3���z����N'�w������%���HX�
���>d�L��0���I)q�i�p	9�� �v|d���E�������(	wю�[�B�8s,!�]GJ��������Y[��ʁd�0����T	�%�1p��;�ͣS[o�!��b�'����PŰQAl�`� ��|����QJ{���H�}�?2Re�Q╓^�!)����&g'����NB��ZX�*�,�s�\�V�!�r;ok[��p%	�R�),�	R Ԙ1G�hO�`m�����Yi�+�7�'so�C�#�8����n���>H�񴁖���HJ9AG�w��Ľ:B�!�V��`�q��?>/pI��yU����ϯ!2�K2�� �Z�aC�AT �x���1^��������ɿ;o4��I�g��R�@�6%D��.��~^��>CjԈ�{b
���!�3�)���/����*�1�<2�)���{��P����
o��w�BE�j�N=�N�ilM!�+��}�SRC0������ׅWemS/��ěcp��TO(���gQ��A�ʏo�+ "��'m�g��.�S@���2[w0�3���(�>�HZL����ؙ�hS9v�!B�%�����8����#��뀣4�3rs�#�3y="4�����u���42#�O������J��_��?��K�x�;�xB�7���q�[*m,-��Q\ՠ�_��6]T�$e`��G�˳��|5��ѹ�7��n8 S���O�q�������;إq���'/�_e�a�=��g���}�=�o��myc:�I:,5~�?#��a8ܜ�q���3�����@w��uɽ���^�����Op?����~u���ۣ;�(fX�`�B�� M��3u�:9�S��!�5rX���h����:!�����x$�R�Af���M$*ߘ�� �l��_�R%�����U�[%��6�)��q���mK����f����GƦUN!�:XN�mȵLH�Ml W��Ʃ�R��6�*�MlB���W��/�C��EH��)hc�mq��ׅހȖ�UְO)�z	dL>�B����.q�3��wS��Vl\����N���n$b�$g��%��E�6�����Sh�]V\/1HnD������ �(Oҡ"�ET�_���a��{��"�K�侱�1�v*d�ӂ��Ĩ�x�|���,9M8�.~|#���ۢ�Yg����8w����Б-49�ޥ9�L9K��HO_�e��>"iF$���^��m
T���#�cvyM���6G��ߢ�?��A�|le� X[��(8��e�U���@eeGW��lc�}0@(6U�=je���a���X���sf��t�~���e|(�ί�E�Npv�Z������ѮZ�f��q�T�������v���/
��>�d�'�� F��C~�Ʊ�������O�����:�W7vo��x@�$��	\H��8^`eF���O�"��omէ�St����os"�pɏ��tq��f�-T�f��LX<��W���a�>�0^j��#��ҊƀHn`�M��N�o&|6HBq�H�����}B�Y�د������>쮲ą�d��ͤ>��7�`�b�陹<룍�|�N/kʖJt�v�ʞ�����?c�k�) 0IC��ɆR�W4	L�(}��JQ�t��ﲩ�l��F����81U���/ib��ѳ=��T��4�.Bՠ�6����ll&x�φe�vï��Z;cb>�V�9�v�d����?4�:d����(ݝ��I#��P�&��`���م6��|�TR<Q��n�1z#U}X�)R4!���ō����1��Tc �wuU���6�\ɭ��6qH�m��Q��|r6�����ٯ��V�H��aZ�J�a�����rZ���z-�3��s����	u�@�sQF�O�pu��5��,-���yQ���ӱy��h��VE)/U�V>Lꞣv|c���*J�!&�<���K�,��-H�<�9�)����D���H�f�_���Z���A�1yC�=�C]֔�"����!�7�U���*��Һ�[�2�-��	�?�Q~F����v��7
~A:Z�v"< �B���,��`J�D��f��D H��>x�OJ`>J50���`<�l;6�(����_E�ojK|��6��rӜXo3q��ᚦ�~��Yឿ�(�ui+ɜ�a�H�gp�¼����%[�p���@�8�L:#g�I.O�!��:_. i0E���)��[�y���� a
'ތ麗jcKZrXֺW���;��D��j״B�FozOnÑ(]~����a�~���ec�J:1�G��a�Rچn�]3g��& �b��,����&�-\���=E�6�9 ��9TKOθ(+�1Kc�ko�\~�Dw_lB���=Ujlk-"v���񀉝��B�r4��݀�A]�%]�ܮ�g�N�]�+�Z-T�kd;;�O�0��2,��0r�V	��O��f�r�'Y-DM�h$�$����������+��Wp�Yϐƪ�P�e���Dj���_�X;q�j����S�E\��Y���i�z��8kn��oM��}{׈y�a,� ɝ�0��L�.e�����	H�`9�M�E��ԇ�[�|m�z.��	G�U4�+������Q��,��˜�:|���½S��S|F�����S�����|z`�k�����u�bl�	)��O�����n�%��W�� �Z��9�dTQ�Q�GK]��sq���p�����ݠeiZ�9��w�~��5g�w�mt�Q�Q���$�utܟC<��aXTw�B2��?w<�mT37HМ+9��5��'�t����9�M4rDwC/)�aK���6dIh�^8�(w�n,k��_@����Pp~M1��/�H.?��������9����H{BP�� a>U�JAe���w.Q�s��5�%�4œ�S�7<�R�Noo��6��i�a��"��Y���#��~�M�7)�8��JP�
ߦ�
�s3��_OX�9p[�c��t��N�.{,^P��ϧ��.aȍ��!��I�ڰ�i�V���.�]R���tڝ䠓m�����~���t�~
���Z��H٭����m��s�zT���G������e$w�ڒ�6�*D�E�k���PtQ޽�;5�Y�Z���N��ݬm�2/A�G��k�`��7��ϵ)K!��?�Kq�h@4�NR5�O� �
_���8,A����y���:�(�r.���좝`���3%M�O����`����x��>c^�}��pD�d�f�ԇ
��X�5���"�D+_͔���T(�"_�?O,^����v����`�1Bk������Y8��@��HNl	Q��<����|�o��홉ͮ��{�U��s�A��@h\Ͳ������UO�����&�V�ˑ%k�t�x�3f����9�w,��+?;�؂o����H6u�}'�
�63h�T,�%{&���Z;�_J��h{��
���B�F���Q�^{�L��#��?�p�ҏ�)��<6�9K���W+��O�N�)��/!��Ќ�I>	=0�Lui@����C?�ݴ�YC���/�e����xEB�@*���K�WY�6K�g��&8':VY�Dֽ��p%�.G��n<��z��Iܥ3��>o�<��|��L�Y,_��]p����G_]4@�7�ǌ#l�G���8��,�kxzkP���j<X%E���L�?�)��Q�زsJ��}��j���"��L��q��IUF~@���	QA�6�I&�8F����N��՘�[K	$�Q�^Y�_F�U��`[(ގd���$��m&�R)jf�;�U�;4�P��E&�/��+�Y������:�Y�q����@��Ml-�r�a�W�o2y�9��90��jZ��h�@Ҍ��6�������]o����s&h]� �1<�C��JK��i���I�4uC�ɉB���u���ZM[8�Ud���WG�:�lbױ�� 0U9���eR�h��sh��}�F�2D�B\!���c��jJF斄I�)��Q�8�ǰ@����>�QW�
=� �R��4[Y_j5T<��ƿ� 3���!Eg0��;釨�3ߞ�"�zv>�!��W�0bu:����Uh�;<XX�&�`A÷����.���m,�n!��:y�Y�>�&˜�}�a���Ck�1�FѾüz�7ޝr7��%�cS���V��@������o7<"�EK��m۾kB�����	"�������%��0�`�l���Ѧ���b��xh�(C1�m��x:�Q�Q��bIQ��C K��X�?2w���Q�*�E Y��G�6�h�f��������۱�r�<+E����>Z`�Wr���H����wz�v�2S�Ps�I���Н:h���f�� MN�$G�2D�c�u%��J���S�Y��"^�P�"R��ܩ[m��ڋ���g�9��W�GO�!�@*���������_�~�[N��s���a<�2B9������4�Zn���1q��:� ��~֩�h����D��R��)���QH(�Q؝��M�v�@���aè
I�-Ƙ��#��H���aoC�t��u %Q��Z��<e_�Q�4O�jd��$�\����m�<�aL�*��n�-��m��518�{��%#��8]ZD�H�s,��=��B�z/=���������p���9�N��e,����h��]g�d����)�b��K	>���4y;��:HK��{�	|W���쫮%�錔��P]�X�3ݗw`��}1l5j�O3���IZ+������E�'�K���;ʃO�D%�}z�	� x*{��j���f�Tt�V1�]���:Ժ�q�3	����ى�X���q�ve��UaN*���*2������W+���I���n�1g�u�������h �:�Ӕ[ڬ��Pt"��u������b���c����SZ����09��	4��KUZQ�g��� ����}���yk�y�P����ZB���������e�uݣ U�X14e���~̥;�.�`	����p�~M�Fx&���� �U��ev̜��t֘���:9RG;�rAD+�f�(��rN��/�-*�C"ݳ���3A���	�ΟJ���|��x�K��TC�e��m�s�돤��cQ�m�n5�\�+������1���U:e$�}�ZI���{�>.���F)�?˜o]��Q��`��=��������z8�QB��%q�����P�a��l�Q���Ͳ|�tD��N����y�AD���'���C?�!����j����_����u���x��:�ܲJ��%
��u�"�.^�{Qr�eA}\[=�Z�0�Zw��˂�CtY��=	��&��p���XA��
E���MQ��_�>��8���F1-2��D�%��"�eɮL#��."�Y���!Ù�w8��x?���%n���!�L���V/�h+�������dL�4%��^��*���"P[:E�Pp�	����<O�Φ8��X�B����rARB~ߤEn(K�Pm��kMDM�����]�_��l9ڰu�J���S�8�M��7+���97��)"�T�JV8y��U㏘��&�.�g�ɖ���=?�r�����l��DK ���lq�0p}p�M��x%�@s�Q��v2Q�l���Ѥ_��F��8�k�	�����
j�+���w-<\XBArf��u��d�e<���kǮ�����
ʅ�^�Mur��8�yŶk��x������bO��Z�pv�rsC��{�}��ǙMDg�\ j���8�O/�9���P�^97��3~l�ޞ���;)���P���\R�1b��Ņr����A���7�g���07|wk^^n�֘C�'�Z���%rٿmdﻥ÷4����]I�?����ȡ�����5�P"L:� W��tUy_��Dy�Wu��uP����]��Dk���J�Y��ʬר��C^���Q��^�Kױ�0-�W��z��s�	=�`�CY������'��4�>��g��ba�KZ�'��s�=�E�ϣ�����qMƏ
Ġ��!4#�k��?��9��[�;4G���� {�.�6ۊ�ݯ��y�s��K�!���-[i�[�vw�ߝ*W����7.��/V�"%K�`�\�����WP����M�>�<:^^�D�o��~��<�_N��?3$�֓��ְe�F �	��z�Π�[e�Ǻ(�\c돠�!�љ�7�[��'�H�4X*5��z�>x�j���:���ǕhCeI!��v����j'��*��9��T�	�#�վx���."%�~$�h���Łe��9���!��X���бn/�ɟ�ձ��L�&�,�mTa�sY��.BL.r��/v�N7y��֪��J-+K�I\ް�/U��I
$��WEk9�Q��\>���^��zb�C�̇�+�<@t������Fg���H�`q���!��`j�4q#����'���;�ϧ:z���.���3��G�Qн�J'!�b��e<h>`KM7�������E��o��Ď!�\��̡v�|f�$�ZŔ���L�q40]��>�я{��8�磹��M7ݢe���$C�r��aB8�`�Tx.�	�i�V�8!� 5+<�r�@U�в�^�#$o>%B�CÞ�Y��
�ޖT��_��!�|A��k�S*���Y�[��Q�m:;��"�=o>��E�:��;H[�ا��P�P^�=�u��FN�թن���rm���Lި�LZ>�F��ot��_�Q���A�}g ��H
B�FçM��褸�Ɔ��'M 2�?�2�N�V[�W���b�_�^$H��e
+���Ɠ��JM�_�d� ⠥Y)�"i�Z���6�z�
�/�.A���8$�E�a)�����;Au2_����D�<94���
��h�ҹ�шi2���p�6V[B��g�QK����)�����7��t9Zm�4ޜ����&Xs�bH$�)@ <�/�N7\-�Pĵ�&lS�}x�I���x��ds��K���4'Uc�3�l�$��.t'��{^k�>̹�X��¢%˫���`�L��?A��k���B*ƴ*n����"�6�fB�5r��W��=�۶�w�Ř�E{���¡�f_�k�W���J����sҰ�֓|�$��a���)�ޅ>t��?x��z�����I�oI�x�4L)��ܩ'*#����->c�c .��H�i���T�枙z}@:�t�F�"��K���8f���K��1�6�E�8�i��/4K��I�Jk7��X;��D-�Z�ѹ�� ��@�q��%�7 @_w���� �O�`dG�+����3���8�a	��v���IE��`Ҳ%r,7?&t�4�B[��XyMos�����j�b�v&��_��i�o��ۣr�^5����^�F�sDwp�L�Z�9� ȥ�� ��R.�	�" ��٨�a��|�.�E��+��*������$i�(Wd/HYn���e��hY>\���
ϥ�G_��`	�ߊ�#��8��=�=i%o�%�I��锖�)i!V߈�;5�j0}m�?������a5-�F*wi�J�5zq�u�F�W-i8�,H�wٱ3�!b��U�6�S�2��+��'��;"j���'��j�B����Q{z^��9��O��걦�c�&�7�i��j�ld�����V�����A@��itp
z��;��iqi��C'���kU��|��k�}gO��ؔu�#L��ǅnט��Ć8$���Ϟ�d���A�DSPU���sc��Ӟ�U�������,�4G�H��+�c(+�s�3Db��0��y Ez�0�:�%���Af�/w����.C}Sg��_�[�r�^){��K
*�8}�P*�۪b�W,S,yb�a��qys�����E����
;vӏj�z�s3^�P�(5��5��!@wD$�)h݋�Q�`)��!S !�{���Rp�@f͖�u�n����8�sȃj�:�x����$WV��tֺ�0��R9f2�J�ʵ�<6����dC���dBG\Gl\M�ڱ|������/4�7d�������-����uE�GZC����_щ�ã���G#�8��N/�`��tEoC\� T�fN��dF��)^�ON����y��$x��)P� �O8.>?w��`��%�-G9�&�/Di6��^�b5�g�.��ad�^��s���,J�4�d���-�j\-���/\��Ǧ�G8���n����L�x�eT�8z���*\)<��S��zݰ�����<�O��:�jB�c�[�')��{�S�����s%Nɳ��1(����0���N	�m��웖�R�a$�n�ԝ�h�j����@�]��ѣ�1C�3R8�~� �⒰䀞JG�t�N��{� au�@G���i$0��tá����1�|�	���:��R�#!��x+(�]�b,؇>�)7��I�U�/f�%�f"�Ĥ�C����"�/=1/~!��f�Q�zX�i-�iQw�=v<]65\��-M����3<2~�>B�G:ޟ��p��:�*�%N���|�S�xi��Lc��|S����k��	�4L���G�Iu�5��n��B�LQ�@X�U�#�1�û�e�B}Whx�Q7�WR�Ǝ��K!�~�w3���������� �7o|Fn��3����,a�0�����Æ�m;��Blh'ֹv���\d	Y D�&5�b�� T�$8��b`������N2<a1�N��_ ~��^0�)�����.4�-co/����6[�2��w����o��f����)�I�R���,ٟ� UK�e9@���H�	N-	9�q��r�4���|�C�H�j~��7�e(w(�v��K������*����7���v�^��-��9��U�r|i��P��^����4�Y�M抜��WIF��+�he�����oO5�|�ɍ��&����4��s���,�Q�e_$����!�h��v�e��*/���W�.eN��4g!��rYՍG�5�p�x�Q��
o?���_?W����r�S��H¸U~ s������s��qC���-��kx�->�́W�ͮus��pi��\e�a��O��~�
�S%�>�8b���lcgD~��n����S�L���߈����>�(�q���ᡌS��e�6$�Z\�&�je#l��NpԳ�o���r&�wܑ�� �/8�0�XC{���B�|ƶؠce�J�,E;r�k�j�=x�R���%������!����r�#��{�4}H��'���j�)�'r�׎�^bs���.���DпN�k�x����4�}��O�lX��Qf��{�Q�G�M��1��r�����L�*��q�4 �	��Mj[�a	�6����x�z�Z�o�;}뤴QT]�+0�R]�7�	�MY8Z
U��.^ ���	��,�Y�OK�e�G�r��r���9I?��� ����%�L����=
�b�� ��T��e����A��
%}Y)��@��G����踾�7�׆>ou�E�X)R�M�7w�:����_?{G@�ڃ������ ��{7TqS,Ld��_��X�>^���F%B'v��~j�V��X�d���nCF�@�S�mPZ������b�/��� �׻��
����(�%A=�ߋ�Li	M����+Nﾤ��bFZ$��$H}RA�[ON��3��vI�;o:Q���Ѭ��y'�5!�����MC�giq�+ڰD�-�A�,��E˛��߉�����a�Q$�0QJ�VN�#���x�mQ(��Z5��
�����bW���Z4������YH���S��'6�'�'��\��+��2T6� ���m�p�`�xn}�6���v5³p��w��5�,����1_w��E�goNhE�Bc�����?�H*�Vԛ��IGi���G��B�,^|K� .N���7'
�4��U�l�?���Yѧ,q]K{�0��X��c�ޣ���[�?7{M<֑o_5|Ӻ����6�k��I��aw?�[9A�@��ǎ
kI����	��oǢnY��陣�í)���x|x5GI{и�����M�	{��]�����U6���(�u��h�yF�81\��,W3�Z��ϯ�`���(5@ŀ	ɬWa�����	ߟ�f�%����2�'� �S�����V���
%���kH%��>��vI(g(� :���y�up���FPk$���Ϗ:�����6�C�+v��,�քD{Śb�5��0�mB�{W���R�1~s`�,�m԰$|�x@��2E7� �A�q6x��5y�@Y��+�}�r[ͳR�1-.߸6x�`��40\���{�����c.�5�bl��1���/�Fm���h
�U�&��g������ʼ(^�\/���Q�0J����^�hN?�<aEm���6�	�݃��I��;B�\A�洼��a��:r�ls��`��G)�6�� ����8_��C�r�Gn;��ӲX�n8uu�*�����fϩ�����A�u�@*�6ykm��� E.�)��7��m]ZX3+zu�
]�N*�Ur𣔘2Ji	R`(�IM���	�i /C��2���t^�=��"��[V?&�v�d�^� J���h2H��Қ�$,�o�0H��^t���aJ�U�����2��B�D1-�A�R���F��;��z��JlmصmAf޻ˆ�����!�AC�̅�\�a�̍BD���4n�A�T�c�1�9=g/�=g�iI{�"�7S3d����5,��ϲ�J'n����x��A��Eס���~���j���������q����U�}�pH�� ��3ĹF��xG���L�E׏3������[�'qX�I���6�����nG��8�p ׌I�|�X�ʒ΅ㅧ�c���D~~�u�,���7���ژD�*�	R,���L��m���T�%�7hu���M{=PGh�"�&7o%2�ɹ6�[F��͒�����������c:��5�,;��ˢ�]j@QG��%����I�cl�S*M;?y�#ʹ��X@�ְ��"`	Ij����{������<T�����7�@��7}9��oR��d�o�@D~����ƧSp�%1�������s�>wJ��p���TME�t�տt�]#�W��L��RBC'�L�ҕ��F�w�	�&�v��ch
��~G�x��	�nH�M����U�l�H�T'� \�F�6�"(���5D/�i�ȋR�;�3���l���yO�Fׁ�_k����-��#�D�	O�9�н�l�����+�D��'���RL>Cr��-�d��OҦz̥�;�a-��C�E�������C�[ޓ��CQc_L>��kc�M!0M�I��tj�(�񧍔�\�!�a�ߎ��u:����a�R�9Fe���H��1�<Y(�t�BT�GG�ld���D*i/�(���ډT#I�Q�@��p@�^?%�$>�\�{���+WAn�&F����n�%��;%��Zȉ��l7��(�Y;�h
v���� ���z�GU�,p��Q�7�VM�"J�J]f[r�:1�A����]�>�9K���QiC8�I��\�zS�
]�X����z?���C�,����!b�f�\�K@���ZmL2�.�gТ?(��kU����O�(	����"\Wt�)�#�	�0\�~�Az��ea�V�uy�EcV8�.����X�obܷ�R�;���NrT7��Lj�]��J�Xd_�_-�F�_�_��pi��ZN�w���X3J�A��1�.��8(�o �c�;�8��b����H�q'b��`5���>�7ʹ�s����"/��D�vvm�1��.�_�;?eǀ�e9�#j�(��=j��{x�2G/MÆ%���m2C�=�pG?����UEJ,g:��s�!���"ȧDl�6 d嬳@0��X��&-4T�1T�6"K��CT@{�y*�Ȍ�bY�n�d� ���Z[�rEy�??���3��DN���}�q���J��7D�8_cU�cp>������M�MS�X�U����7��&�:�c��	���Ц���%����Z����K�z���:�B�棫��-ў�x�m�����U
3�q��({��n�ԓ<p * ��4�>��E%����`��ZAF[��^�oZ�  �Q��=�`��4`!�������}��NW����1k�:Tq�J�:i�̶��q�S�-̀7��*�T����OD��4�z��5�c材G�k����_���M����@?[Ih�= ��0�u(S&U�J�̅>L�CD#����q?H���k\�����_>���[P1�B"S*����ֈ��-<�0�����\1C��^ ����-�O���0ײ�֍�)���|v�v]�_�>@F��Ӕd/���\��(���T&sj@V�F�-����� N�ܟպ�GP�5�u9;��{+�q;���G�{�0��PLu��r���\'̐������%l]���V;*�ܩ�9"X:�O�q� ��F���e#Q�[�r�>��Qa-���!X�e�KտYFA3o��d9m#�0�^��
!
ь�+�����uD� �e�xK��B;�bz�@"�e�)y�)�b2o�z&_�m6c��Q�Ց�����������aL��`��,�Υ���Ę��6&h�����Ժ��p�{4�̾}�`4F�џ#pR���B�?����Jܾ|Е�i7��� /�219��L���<<�����!�"J�O�j��Nl���>�a�����$��*��y�U�P�L��m�{H��l(ɎUK4΢��7�sxz�S���1�-~��B�[M�jLIW�݇��ȍ�R�ά��I���*w�rKZ��8���\����� ��
�T�!�֑���E�^��zN�ژ��c|�~��>�i5�3	��sϤ�G�4�/1���]���_�'�k޵Y���g%�y��PB�_�Ǉ�8�ԥCmY��.���\��`��������(I=�^�Xr34�I#ZK��J�����eĮ�N�d�i��!<$���>I�8+[>C+1�7�Lc1�=Y	��p5m�5[���Uxs4A��)x�*)�~�]�������A�M����,f�*8��U}Vm�	D��+=����j���ݕ&���XQ{Ѓ�[�)�����e~ os[����������S���y5��V�Q���^��!��H�!Z{���iC��$Oєx"�z�b6�me�p�,A�~�� >�d��r8���i�z�}��<���g�5)�V��;A>��.��C��T-z�3f8����iU�!�����![�T���!�%��C�c����>�{	�բ�OMp�?�+�g?!���/��I��S.�拏�C�NN��/�KH&��$�/��p��M��]��u8�-
T�rH���t/\����GJ7Q�Y���'E:j�bq���_Ei1-����_��:��_ƻ�]�Pm�+���N(7[�~R��EK�S�r�/��\^6��Vb}mW�C�Y��G���\{)]����ѿQ&�ʹ�N�+��7BU �`v�qћ�k`�%T]o�P�E�,K��5U	�H��t���@x�M-h �k\ZQi
q�f���Ӛ����S9��S,��^�1>.�{�'���0P��R,�[Z0�xy»6��jS4���!h��	 kR����ӹ^�Fj�OB�eI�#��l�h/S�� ����u���-gN�b�ƛs�!���w O�a56Q���H�?�F��՘Fe� w�Z�[����E��# ,����1���ϥot�dv[�����D��p��g���!{��(��ʏJV�Ws��b�z�<(�-Fe+4S���R���X��j�w_�dV�`�n��̂�X�uY�a\��U�i<ʇ[���Y3%Ėi�q���o��|rb��)�8�_��J�R�F��}+��t[�[8�wb�4"g��ف�M�4�;����TF�;L�T���y���Խ��;������ʱ��ϗ��y'�*�$K��-e��@���HK�+V��'m����Dz���b'l��YuvF�5��N�c��WkTX?���ij
��]x��&*���x��t��`�/���*̖�xS@*�>����+�J�m���?�,'�����i&t��"�Oe�Gynt�Dѹ/R�_�M��F���Y
scJ;�!���L*u���%fď߀;��$���+�7z8�|�=S)��;�9Tj-�`��:xq�8��u�sb�Q�L�"���܎��M�O#������y���qI_/�u�J�Gt�Ѩ��|�:L|�H��6	�t0�.�l�g-�w�^i+}����Q�nl?�V��.�W��v����̨�8�$�`�wg������ߕ������ɺ�.��&�m���%\Q�:;>�
H�}�F'�e������%VV�b�d���UxG����Y�7����"��vɒ�U��X�����5��=���װ�E٭ /C�Nd��xoKϔ�>hH�yCbP��a�x���6��j�\��3J�h ���� �*�C��^�[$��og�i���!�a�5���#��hN�;{����6�V���r�NZT�.��if�7jN����,�m� �L�RU�������9n�]��Z<"�j݀X���]� 	���;6 �0?�u*��)��s�l�?Η�: � [��~����S�'�M1�!�[Mw�,^myL��z�)�<���{;��؝dz�<��:���M��$
 nx#�X0ԷUf� �?D%G/��6s#�5+A�"���g�	j�I���`Τ"�3���x���[���_"YN���wˀPSG;����q�(�!V\j�=A�W���o�vs�v^\}�2����͢Ar'�6W35T���SZ��'j6V�~S������%5Oz�J;)��X�
,f���۾p��V��P��8��`�	}r�w�b��ǧ����
��7ڴ�����Н�e����te!:�ʤ"]p����󃢠Ϙ�S��.����XL�S:���|��Q���2�Nop���ĆY��e5aFA.X�����7�T�g5�ߎ�,�E��ea�C��%��~'ވ��~g��vn	���e��J��HY>�>H�௷<��ԭ����i��r����ҥS3#_��t��욚Y!�T&P��?5��_�|��:SQ�i'%$�	A�p�kU=�>M'�Ԟ�t}�������.Wbk�����YC% ِz�����T�����9�P�j���k�y�n�Fߤ�i)���o��=��:���h�o����H
b�(�8��(Ѕ�fZv[���tr�aTkL��Օ���7^G���zm���n�u7��e��l$L�ki�y���T��B�u�S�Q�hXM��_���mt�+���C�Lo�O$��\�:���^�P[�j�H)XL>5l�Z{�&��hd��p�^|)a�6  ҚL*�oMC�5���?=^Vaw���l��J>�
�!��� L�m����a��~�%CY<�0�˰�SK:+���ߐ9,�Kj��4�
�	t�-V��L�'C���2�W�?��Sѡ�n.���p��&�+���@�wb�����+�C�;����t�0"�Y�1�_e�����\B�a�%���2�FB�h�1�S��������V5<��f�X�x@�g��V)��+���l[��]n��R�ߘ˼x��RmU@����uO.X������2'�d�������(A�ȸrO �^��x���.�s�ܻ�wC�l�Y���h�������МcC�Kb�㹟x2_���5�Cc��)ضdVk�V%���oÿ�7r@-����;�(��(�3��\Ye?$�75�n�/��m �&�xa_6�_^I-@n�����el��(�!✦mM�B�3�I�Ӭ����)�:Ԟ}���f@� ��u��ˋ�W�~�5���3�^�r!~�z����$��ĳ�C9�z۰�lNB��p N�j�F�
p�x�U�+��)K��4;�bK(&���Ƅ�1ş?�
��"���n&�P�4J�}ǲ�TV��^KI>���)=��<�^' |#I 2�Ac�Q��v,�4���;+�{�2����-�d����f�R}0J���28�#�Uqg��m,k���d���H��JT�q1a�|i�k Ӫ{^2	���G_�ު$%��O���}��gmNG�����|�� H�D"�?�<�2��r��~˰�:kc����g�X�Z�n2�� @���>7�/���.`(�Ze8����_���h�w��	7�=�X�Qe�_��H��"O ��Ґ
=�&-�RU�o
fc�W=���$�>���@u�%�}mHY:H0�(�ͮj����ڟ�ٹ,��
��J��m[�n��Ky���m�	�,�a�W�~�}P����NhG��n]CN�3����(����'m)��MG��a=�JG�d��ЪF\Kt�Ds6���ll�0U��r��+}��3�i�l/��/�˱@"������>�L-��ow�3�Sy�x���������Q��q�`��582�O9N�m���A�����3Q��V`����b�v�~b��4������ ��	%�lB�H��Г^v�aB{#0BC�v�(:�����1�h�� �[�2S�Xda�u*��D�cW}ߛı,dM?�����4#_I���M��n��[�iڃ2�N�FV��Pض���������E2+ʜ���L��1a���˅�/h�`B&03���b.|��&Enh4O�������`0a^/빚�2�VOj���0?j8B�K�B�o�q7FwP=#��otN{oЫ�7D�ѵ��u4/�����$��F�'څ�G��,yz�T_����P$0U��I"�Q��-���{N  5��~��E�' �`�#>��a&��mu��z�k��3�n咹��v��U4R<��űC�LV�-�F�I�i�����G�u��w�#g����/~:��V�:Y��Æ'�ݪ#|����4Ng�v#<xO˴��gE�S��D��/K�6$����[+�v���E��u���'p� ��d d+u�a��߭�l�Nz���ًE�.�������YJ|u�1]��3��y�⬟��k��<y����{I����+���䞹bHņ��.�
�gtm؉��N'�ol|Pnm]�E�'-���:ͨ{@��$�������T#��������'\�V@㛉��ɦ�t<M��녟�����$���pӴ��o�E�����>:q�)v�1V�UK�f���-tp��V:ns��V�&hF[�5�=c}��Tr��RV��B�������^I*�D'�'͚��"b|0�'ӄ�
��n���ܗ��JU\��HV��K�h��ͱ|'$hOԮ:""�S��k}͎�/'��)?h�Dz�AL���k38M�P��&��3$Ta���}�O���Z{�i ���l�{�K�)	��g����CtO��Q*���v4��OdR������	)�#6��,­j����iT��^��j[���f\�!�3��o��,9%T�PO5���z���ĕ�t��`x	Phi"4�j	�S��D�&�9����K��������_*�鉔�z-��^S�x�.<�����M �q~ւ��l8ŗ� �lo���p���������X�놠��hN�(ʱ�9�9�	QG3\��fF�,G��Jx���T��P=�$�����t����d@D>P�e+��u ��V�k����C֠���q �&PB/���7�Q؁��L}FtKXC�7����]����7�B6����aZރ�.g��顼60QZ�b��Z��r��Ѓ=��_4�&1Z��$�;^���Lq��Y��]�.�A5_�[�-.�ܞ�!��X��>z[��1��686.zM v��j�Ϫ&'Gܚ`�7T {?m�L���_k�r�,��T{гeJJ�y������]����b��Q^G���P ����W4�v��ʥ���0�\2fy&�+�O�p<��I� 2P���۠lG Jt�n��B�� ���VҔ�������c�k˭���(�L�����@/AY���� �k��#P���z�ݻ:�-��3ޮ�ط%	Cg˳,Y��8��u�&{6=�s�np� ]P	�=�>	9�8�%4`稍�f��	��
�(���l8�7;���ӭ��lD�xx���e��2�_"R�2��?�����;-3�n�������+�����|�5AД��J������6s��v�~�Օ�|1�4��ƌ��_f��B��e���Ԉw��}��1�pFDz��/	�����oJҳL��0��H~Ӷ��@��{�1�r�DE�oʅ��sH�{"u�����^3��\><����/=S�+��8����9񏢘�����[�8��휝���ʖ<.xm�_�s�ލ"�D_9d��5���}^X�<� W�R+��Dã��mg��L�m�;ו#�D�2T��҂�o���E�p�YkEWZ���%���wB	4 Ua������]�5�\~�v��D�ݢ�V�#g�]�!B�*�����4��s�T�Bb��4�v~x�F񙡾�`2�}i��A<���o���k4j�gGWN���9��Q��^Md�G�����N}�j=���ٸ�
/������r�*d�#-����I��%�\�z��0�3���ر�J�7뼿�R�7j���~Px@��u�
�tZ�Ҩk~, �Oixo��C����EO���0��}lt��%(/m_��z�Gz.VYY@W(s������ �{	��)H�v�D��\��\��w���g��F�I���R���;��}��u�o\:aP�$�B3ɃJ�r��ge5�lT4r�_�AKq�خR���JD'�L�AW���o@kL1�D�\H�`n�O#�e柡����Szcte%�>!$�o��yq�@�Y���!l��c�(��M��O+G?H�He����4c���)q[��R�)e>^`o
�c��� ���]�O�4�PE�BS|s�:��-�'�q��ԍ7f� H:X0p	�\�d	����S�1'�TZ{����⯳����!zyR��17�G���-���������o��&k������:��۲MD[�X��!�7�p�uq�uht��X�A����[�\�Z�(�v"��V���ʏO}�3�B/`pg4�X	48�Xq���Y��'�K�f�%�?�(��Bp������&g1�O)��A�����c+��C�5�����U���� l�S�})�Ѳº���̬e#I���ðN�R^Y���N��(������>��O��1�4�V�)��p��{�<5B�{?��
��(��ģI�+2�'2V^��;�f4c?P�#�	���G��,�ے��܀���'�#��z����u�"^�Wa6�g���F/�:���_��x3	���+�w|�;�dصӬ��Q����a��xj1���P��mn�qS@�u�ֱ^�5t١]�8��J�&1�"�~��x�.&�f��3�;���ĸ��%����D�����#`:H�����4a�1�CdeD�m��}޴���!ztb}�k�!Z�"��J�T?��ߴW��9w���Yd��9�C���#�����c���ZN��.���5;G˛g���1�+b|]Qj���� ����o�U	��t�٨�����Ȥz@�ۍB�~�AN�aH�h�MA������/�؁���Z�
J�
�h��KB���]��ȴ�ì�M_�)�L�.�V���:��4h�}p�s��n��@p�΃���9��|=l��q��͇���H��}�쥑KXd����Y��>�!պ�XMI�^1i��u
�J��DR@d]>º�G6�Ur�e�	�5<�)��]�.�	{���r���m�/���J>�F�:Р��@[�S��Q��j{�ߟ��E�P�7z�>�Lu�\����S��T��R��
�)$��޵S%�K(ܭ,�5��c�G��֥W(:�,���p���8 ��Q�MNd��W� �JFb��KtM��v���G��U��0>@���q��<%�)���t+��T�f=4�F��G�0��Ns�^�u�_�luś�j��Ţ�*c%V=�;ǴIN�����<�֭�,�n/��X>�
�7X%�wǊ����bM��& v尀f^ѓf�Z��]$KS�hX@V���E�
��� �s0��, [���I�Ǝf��{=�a�zw�e(U7�6a	�P���z����k�O�U#$���  .)��U%S_r�����T�>�=��N~�Rg�9��d�"��->ȻS��;8J�D(&׏ŋ����e�yeiN<�S:(��l
���<)h�q�]����0zP�f�t�1�ۂ��7���r�7q�H 3w^@/�c��wpQA�`|�@��Ɉ#��Q��J;ٛ�:o8���(��%qjL�|>GW[�ʭR���d���=�1��'q�Hݡs�������c;?X�dA�^ ��W��b.S�wI%HV�p4�~}�.K���|�w�֫�QB�{8�;e�R��[a%05��_�xG@|�7�ndw������!��a�4��lAO�?]���J�5*��SϴѼp˧�O� C��fN��[*�D�w���O��T�\�py2�sة��	��p�~��Ag'�� �x4�M�l!���W��ح@���bvi�$@�8f^N�T$A )�!�4�F�f���E��`%����k�p�GJˋ�s��d�{!��d#�@��K�����`#�d�j�����%$I\�W�����:^��|
�vȍ�:Qu;ZB�qe�m��C\�0��G�H��Q,Jf�A�ݵմ�����eXȭ29�6h��Î���h��0AM�p�!�B��J�f���*\�)֜Q��Y�h�=�b��+)AE\����� 	��76�-�^#�=���VK�E
�6����I� ��x���KTPG2MЭD�k5Y�H�B�e밚4sE^ �$�ȉ��1������[v����zL��#MJ7�V4>S"�i�܇�=����$��.cQ����g 9t�����1��I8u=+�x�:�q5Ji���<zI���nr0Y�$2�����LU=V�[��pLZ&�*�g���~z����fm#ӂ���6v8V���n�I��\6�W�.┉�y1�j��o�LG�ݘ6I�e-�YU}[��#��/���MzVYZQX���ĸa�IDw1�xC��UM���\�.�ۋtb�1��w�UmMuh�F�&�b��F�	�V���L����x���)iu��{�x��/`G �z�T8���I&"F���A�`|1�(Msk�ك��I���͖'V�N�*2 }Fa�e�!�� �(� �!��5�Y9��#=K)=h2�Ԏ[D_~��#�S��ٍ_ۥ�gTE��(:
5��Qu<�TB�U!+���7�����ɫ�����c0z���{�ta\�F;E��"�6c���L|<��������,�};�u-�mJdJ������zԼA�����j����9%�V<(t4)�T����} ,Sӑ��9�M%��s��<Y�1C����e�٢�H���J斿z���ت�6&�/QP8VM�7=�!a�UJK��N��ǸX������_.���(�{�i������3�ێ8���h��15�l��h��;��x:���H*ݱ����a�E���=��8I�;3���9z�����;iȗ��Rd1���$j!��� �pqˡ��0$X�h<�1���gF����!���_fB�2�uO�:M�ع�gB6�4�E�`웑��ɖ�5�J͚t������0�������`�%;HN8����-�]k���M:�&N��UjO��[� 	��.x-Q�r.�eQb;����Y寛���� )�o������,�fn3�M|[a��jA��u�֎�+ �4��f{L;�e�Y��@�W
ñ����f2q�U���t�y�`_H�.��jn��	�TsQ;ua���s0�eb��f��s<x�#�k@2 æ�'�
t&02�/�' ������	�,�s�7Æ�S/��{{����N���'A���S$h�L����B�����3��[Ж(�=*x�e�FhOq��-������?a�>`����D!�^l�Q��F�5�,:܎'Ӛ1���}65��X�}��gP��ĀF�~�
Mvt@�٭|�&5U�02W�RD-O��Gn+��;.U��R����ʚ`���k�$���3�īi��خlAEb���i�	��ּ=�49���z#^c�ŁX��[��d����MkK�Hƕ:��{�X?J7J�Z�*E_��k����Ps,�	Ǹ�֋c�>	��s���X���}��[��Q�*(ږT����x��F�s"���Zz��+���f�����l#R���Gx�y��-�Jw�ɉ���5B��e٢vqb�h�9@|C�#��z�D��&�O��3_�\�oc�̜u�9p'�#������]�V�a����JmM�n	�,C��Zc�f�$�&�/��#?�o����8`n&����k[g�&�Q� f"�7��k��,�{I��ɯ�Y�&��G��	�a�w[+���ӛ���F��=�j���������f�f/�3F#��Օ����~Kـ�O�'�ׅ��Ph� �\��&-7`��Y��R�K��U�������)1�W��`�F��x��i3�n�+�0G@��e��ߐ�h;�Q0����ᘰ���>q$*����+��D`V� ��ШF��|��S�ɚ����Y�9��w
XHCw}O�I##C��g>�E(Gg S��%�E�M6�ٶ��u?�`
�7J5a�)���ȷ� ��p��qt�d�E���!2\3���a��O3�2���J�;	���\�t"=�[]=ఖ��c�p�\��A�,�,���Rn�X���
�x�"�zcٓ�����]pI��zϱU���QW+��DuxwҪ�0Q3�T��%4��;�Z7��{�)Qb�ze#���qNO�[Qw�M�x�L5���%�G�ڢ�KӖ}�g9vGݰXn�N����ToCL���Z��M�I'
»^�I.�"%���]jJ�h[Y{@A��o*:��<�^<��u8����6
�7��<�nI#*��&�����{�u�A�?x���z��@,�Ɛ��ᩉL�N�=T>��E������y�$������*�e�I=r=�IÓ-�7/���*�>�rz�쓬�����o�Dl�]� `^:l��q��wM�*C=��ݬ]���I��[	�J-�uv��-�a� �dk�����JN��i�l�Pv,�b�4=H��f~�p
L!��^!l��$Q�$o;.��!��aЅ�/H��^�ޕ�d��)p�0Dm�J����j!��;q� �:�>�� �v��1ØY��܈}��[%�m���\���m,�������=F���7ܪ��N}��� 7���y�{ADId[�2p�t��C����%'g)��Ík�.G��!�ܪ���|ג�Ck�͗w������<c�{p<y"]c���>ӵÀ三�zV�9lpz"�Tl�!�z� rԲO�
a&�
����3��]�}♢�+T+	rDN�rQ��u4E+�r2UIb�W�5�����A�p�쌗b��@���Ͷ�~��a���X�u�a^�u�I�P�m���CU�j]cfμ�wل"�f��R���뗽W��:�X����y9���:�V�D�������kߦ��PuK��b �����b'sa�U��8�NL �B�I�i���_�r�Jkh1:j�B�U�ƛby�K~����B�9�[��w�С���Ee������
ް�u����)��Z|+�L�:����mƮ�C�@�����Qϔ��s�o��%��;,��aRg�z%�n�O��Jy>�>9�e����f}��,D+=��\�N�a�f�f]`���
6��A�Ru�Vi��]g��R�X<�:���Fu��R��vǅ�l#�ߙ�	�x���#��qoDN���#��w�)��8�=�����j��K��&��ՅXz�jY]5���p����ty���k�&|�{r��gGED%�u	�pQ	W1xU8��yV�=�����F'F�o���Yp$;����Қ�l���(i.��������a&���8�P��hs�w�co ��-��Κ�)Ŵ�C�A�;�#,�C�g$A�_�����L[+�	7(�hc��TUn����M,�h��ׄWϕ���XV���2?�Z�/4{�Xh/uCn[���;�������s���mc8�m����<���]f�ԣ?��V����Lp�~���gC9�h��V�O���w9�rM9�d���� X˙�f����8��b�rb<N[q��Q�Ш:SE:g��s6�O�r^�£�#�0F�[�;�;b'�&_vN��SzM��Y6��kJ5�oi�0��}�8g5 ��ڢ�]��}������`��k�#��D��;��c�h��e㶩�>�tc�jٔ�1E.-5��<ȃE	�иG_5_������O�YeX$Ԟ8��PX�X�
y8��ҽ�״�7�d�81���4�B0�k���cR4�"R��RRz�t�����^�X�5��*�����\Jd�U7o8�������1��ͺiQ5rgY�l�� ���~K20m�=<��w�,�p�}�MiRnS��.5��G�D
̃�n�޶8踰����t��q����[U�C��1:�x-G?�鱰�5gpO�Ϋl�b���m�/�b�jR��`4C</�=EI��i��dC�o0�W�5uY�Ci.��.#>��b��� ���鮦u�p@TP��d����R���U�zb�/��	��2o4�1ҷ%�$�o�p�4��B���E|!��Œ��GF�Hl�4Utܹj:Cr%h��`1�f�����L��ʱ�0.;��k��kD�P$��5Q���V|f�%��`z ?��!1|������k��ǥ<ܘ3����b2�꼶Ρ�d�4��,}���O�ϭ���G�'���.>e�Z'��~�p_L��݂�z������w��&F9����-��Hl)k�ܾ�d��^�w����I�S`ћ�B&2�Ya4������lo�_��h^�r�$ �8� ��}�>$�x�hs
��z��p�s�e��Rݣ���n�Ꮂ��C�����?8��{|	@R�5�,�|0�tO]�qef��z�s���O�D��1@��X���-�9�fm��?�ϻ�u���2#�Np�i/���a�+[�f0��W1q�e"}������4\;��N6�/��c���)���>u�}!Cp96�������-v �I�K��^�	սLg��b����􅛩��[�CZWΤ첰 ��đgU\�q���1I)(lM@Q� � ���u��U+(��������%ڏ�9h�P�A�m�o	��Տ\m>?�ϙ-fx��j1ʣ)�ޓy���$u\�0;����9O �r����
/��VH�Q�hʕ�3��qU�֦���^���~\y��ʹ#��}�/''L�g�؇V�����9@g_7<\�N��;T�bv
W��t	xј;�V΃���pP���uc�6r�B�9x�*#>�Of�f�2�J�����+\0ƥ�����K2UH�&�&kǲL �cX�����׽��8���������#~qoq���iֵ��2 �2�i��v��QI�{���k�J��.g6�nc��u�I��eg�0���MV.���Uy�J���}C䶡0�`��ӳ��=rdZTH��[�ͼ֩�V�j�)ô�>
�_�{-G�Z��[��Y�uo�槪q�W���Hޜ�yYG��*h�_�b�2F װ���L��h�v��7�#g-�-�ۨm((�<*�+�b����_-���{UmM0�>j�_f��NF�(SjG.����4�O|��H�I�\�#�ȋ&(��+!�p���H���h �ǖ�oN��B�x���S��3���+�.�}s�R����Vv��t��>��0E'����]���^���4=Ы)\���b �{9�����i��ḭ��+X�.����`�a����#ҧcno��t{�*�Wu$"��k��`������v�6]�R#���w���vr��[�$�Q��(^S�u����x[���fDY�R.�uc�|o�'}+�f� �|S�#�2�w�"E��}���5Qqu�-Q�5ƽ\�&uݫ�&���EB��NS>/h+-�e��;�3���p�2��eX��L��0\��"j
��{s?W�RH�LӢ[� �U�g��'���Y"j��'�oF̩39j�0�P�#�ڊ+�"����~��E{�4=Ϩ�jW�#bD��M͛*�j*���c춋����A���T��(cbլW��#�w�l��W7�m,ئ\X9#W�&G���>'�G{����k�	���y�䕅M �|SR05��"]���}�o_{+g���>}��?]�ʷ(#��-��-���`��w��G��x���U9�]�~h/b��%u��[���!'t�e�p�{�v�&}7�����O�P߁�=w�F\��4�ϻD�5h������W~J�.~���?���x� �6"\<_��i�Z��"~�Ο_S�%	^���(�Z�-�u�	ſ��Mhwq��SUnݏՒ�б��S*p ;?4��RN*ӘR���f����:A��;���<�88Mik1�V�C>4��2,8�|&�������fpJ =2O,q������^�x~�hf˱1���V�Ӿ����J�/�A:F8Z++����6R��dL�Js���}R��]�gJR�M�v���[�Βk�8�R��0d}�2̻侣k&�L��G�wq��!����-�a�f�3u��y���ѱ��"�>:.���qn}$��Y��������V�=���<!�'M+O�q/�Ǩy��B��&�"�b�\�'��H�( �¤��p��e�,��1� /����f����ą]sd�_[d+l%2%$�}���S %����r�h�+F��4^f�UZ����Q1�x� ��\�{�>�H�D*6�ټ7.�����-�xU�� ��M�|�A�XB#iRb5�Ĉ
��4�;�8h�N~�H���;S%3���f,�z�4��f��ՅZ[o����c�f�2�)���Oq�K��@��Q�zl��6��� *�y���v͍K�f��X!5� Ԝ��n~b�C��6�ߢ3�p�V�W��pJ��t�6�%�/n��n9�1a1���@G���M��<�?Op��2S���ә,Dr���خ��6�χО���2�Qo��E�2`E�K(�I�&�-�����T��	�
�}�C�Aw�;�,�˸���ׄw�!�E�R$��̒��U$�����Bl�y��L���!X/��!5�Ǻ��a����C�䟿:���
C Q�[�x��r�{�`�d�s�?�15E�d�(Ll��j�Ƀ�/����ƀ,�>��z@Q�D�۱���K��#�j{��Mע ��^��`j6�@2�������ֆ�c�\��~0��μ��އ����G\좤��K���	u֗�{rj@�_�'�b
��.q�*�x�\��d��#�u�^�z�C|�X_ep����5�!���#`FX�ϩ�Vg��F৬�勼���[.�us�ㄏ��2`[PF�Qf5h�%�����������>=���A�VxƖ{��@ �c,�溷��}�Y����g�Y�z7��y��eT�g1gg���-��gi�:�j_�/�Nz�=*~&��/�4�QϛO��@�۾ �j�p�'c/)F��
z.�{-'G`�����;F��)=�Uț�~yg��f����^%V�O�̩��B�Zz�|��r3��Wod12�(�@$�uy���-�걶x�t��[�_Q�uv�L��\���rU�P.��l����XRS�3&Em.�f��oӝ���2�������٠f١�D5��
4�˽}��-($`V�8� !�#^L��Ü���(䮰�Զ���rE�]�i:H5۝ݱ�FU�&��K7��|3�ܧ����G�L����;T��;��"\l�z�� �﹨�y��@F+����3A���Fݯ�j���-:2��8�5F�چvm�L���Fھ�C~���2�d��
y������l���H�S�%."�ZD��B)�������e2ھˬ��mo�yEg�GH�N�,|P>�t'�zZCS$nJt��]\���xt;�`�xW,��WP�N��ڤ<J��pu��Z��$�Ml�����BF����2b������)L�ڿj��<��ڹk+�$>G�()��O�m������Kz��◶��������ax��R��J��p���ㇶeϭ�\֐�
)ȫΥ=O>��;�dx���6�ȯ۠��m�}&0�>)x�g�Y�A�3�PRpBK:b8l/[�Jhzߩ�T<��c4z� �;�ϧ����a���u�ڍ���~7���Sr��8���(8�%�G��!C*SAլ2�T��S�����e���NO��+���J��2`���yt	��kd�	�D���u]�t�TvI��D�m)?�⧊f�*{����'�a�S�L��C�C�ʻId�	��+�sZ�i��ԯ���Dlr߸���7ߌ|' !��0�$�F?���>��9�.0�[|QQ� و�YM2�i'�붴��Vo����O�Jt���Z�[N�4 h���h%NT~��x�꩎�s�bV#�}%�|���T��lmT.�cx3��C=��k�CdYa+��6[t������pq
�������^ޖP�8j�E�Bʖƶ _���%is���W��l���;?��x��-�ރ8U�Ɏ6
��{|�p6,����@i�55�_�~ ��(����a���Փ���u% ­�ϓ�z)P�ژ5j����ޔ�	�ʼG��A��IR�efiޫ��,��(x�����vcyć�DQ���tl+������4!7@<V⥂�M������V ���}�������Y01����]���D�{VN��`fh�M�\;�M��Fd�Y���Џ���)��z����èa�y*~j����f��M-(��N�����a5�����jT�7�`)������\��պ=6/2[(�wy���O(lC�f�M���&��������w� �1/u�h��]SA!_��u)�c]0U~shS[�!uf�W�J0��B�.��P�,��7�5��f�c��t����Y��/QԴ�s'�G[w*��m��q�	�ׁ��7&��D���U��f	�}��{�s��U�������;ʗ�}�� ~c�Y�������v<�E��T[���a�(86 H����������w%�#�hl�@)xX]��sU`+���pG|l�
�QX��x=�
��r{���i��n	�s� *9�Q��RƟ������H��.8�*i)��D�p]2E���G.ۗ�q����MU�CNc. 񎛙Q��$u%	�pE2푢��������>��Q}$�	�W�g��o��� �j�t�����s'qV@�h��g�>a7��~��ux��w�o�=�[��96����+��ﾨ5�f�f/��]lE�=������7���\z�/aR`�f�����g���.��S ͉]_FMn�F�Jg��Vy7S1� ����@ _M���� ͙��o�@���$�i�k�u���~Jp�&E]6	;]$kH�P�[��H��	0p�NR��ܬӻ	/��v�����z<5�ç.1�W�ߊn�6����[�%$ �lLȉe�2V\9���y��m�5_�i�{�Rn�Y��Շ��5�O�<~�$7�j��K#K�>^�����|�	���`"e�Z�L��ewk��'~0W���0L}�JNH	I��{ML�Fֵ�J����
qD��^��N$>|f�J��&�.�p�,(0��\��3�u�j7�_Kr��,��ҙ0]Q��f�V�Ӄ��r��HӜ��L'L�[�l("�e��[�I��ZvKSPf���C��,������	#`~|�y�iZo�r�UU-&_6@A,x[��/bᇖ� pE�:hPos�I��k�26^o�I�w�b���&�@���S�_xx�kgܴ�Ly��P��*UXa-��ɾ�!W���D���a� ��陀-�J�U��V�B�b�<��d-�Klg�*b�<B!���p&�1��I�ʁyY!��{����u�7��7��'�c�r����SD/+9{����6�)�yJW0�_�l$�^�ER*�IF\��Nd����@���.]iB�Ѱ���A�X�wE�t-�j>��Ä�x*l�߫��s� ���,��3�����#�r�>=� ѩz:T��'�
����9�	�ON����|Aݫ́�0Ы�4-J@��]���n��I,inUC<1$����H�IG��U��	KLU>u9=�5���|�
KLș�Y(�KVD0,m��8J�����#����VD�K����+h�=�>��a�Z��$=&e��13�mx���߯��jF6K���U�8�ʔ&�g%�Mo<������X����������m�O͈6}�����1��%��x��p�m�O�^��Z��9�^�"Ѻ���Jm+x�J:�oB~� ϿP��Zp9/mf�7E�c�(#���Ov�=y�%:�#�y���#v�UT�MDȀ}
�0�n��T�c�VF���������x��d+K��s9�Q��}�(�/6�No�T���3^���%�b��1R�OVN=4�]��@#��&&k�	R3�~�R�n3��V���qR�4�}���i8㈛�z�quD�#7�z�9i�v�Tk�4 3��iY3�喯̍�%#�!�'IF�\����K��%�Kp��(�a&�Z<���I5��h�E>Eu��R��o(yC'{;s�ˌ��r�����6~&�Q6�T���&�� �� ���xs�yB�PRno�����yAТ�:�\�Z$˺P��`����\��fj�P��J�Q��Z���HQgj�MO�U\��tw���;W�[QM�� r6f��|�@�?��I�������T��ݾ>"�Z�Ly^��;l̈́�2�Șъ�����T��.��(E#�� �L�a��f�����q�2�i�a)�ĕ�s9E�;�C�����_�cp��e��XH�s�b���ZUf��ϵ�Y��S��U@j�_0��|Z*�
i\����u,��
��#�:��y@D���9�,��RB)ynVB� Y���Y��e&F�mhUH��;�=ô�4�����uӌ�
��`@z�������C�0��xhM�a���S����dL�,(�q�vaZ���V����l2��x�= k�Vo�t�=<��u�Ǒ���k�nr�6V�^�j���L!}�����jމ��������wx�a?@��k����
���5G��[[S2l�;f��~v�l	qo1�����`��1��H΢��
[�ym(��0ݠ�͐-�  �T�#.��a���ݭLȖ:����'}�ҫRs�s�(gj���n�y�Э'�1-L��Ȯ֬<7۷��������2�~�qEl�BK���vc+�tC�=�4j��{UZ��*����/�ȵK��oͭ+���J�g��H^�L�G��) ��م:�Б��?����/��:[��}���cX��@��1���^O��͓�f�*T3yj�����BC���be�ԝ9h��|���C0��о���������h��gF_�aB�s<!��~����Jh���F�^)�UO�)X"�����'�L8�����첰��O�&��j�{y�<#ƹ�)�:P�1.�1��>V���$
f2!�9�Wl�X��ZX�w���̅���YGLY|�PmS�l*���2a% G�U�yؓc%���闬��KH���cM�1��t�����O���s�����N5�Ĉ��������c�/��sѱ��\ąp��S�6_�2��F�p�\[L��ﴐV3�r�)��4�m����o���M�&cV@j�g9�k�A%��ȫ֟%#>Y��ܧ/�w�1z�ޗ�2�<�f��3]W� ]�����T��w���C���-�\����"���рi�qm�	ďϕ&�LY�|�+��A�_׈���1�p�o�\��Hq�a��=RYl/)ba�{������Df��3�m�Ш4�����(�=1�ԳNd��?;���,&G���:��ʍ�{������n�����3���x��mD�p�L�P�_C�\�P�Q\%�D&-�R�j�
�;��8g�8�>NMn-�$����Q<�����B΍~����g{d�� $�Ӗ��(r��u����}n��;�A*8e�4�Y�:�Y=*|������[7���kpbY{A6�:[��E�w��z]�,É@�W�%��Ӵ6p�*�͒T���Mfi����w!B<c�m%u�/O�<�u�c���W�E��l�xX��!��3��XR�a���R#Lh�poP�WD�.M����^)��:ؔ��T�U)y��V;�h�u��>���3���*N�uQФ�M�u�j�^B�y.�b����}j�V�����I��ߵ��L��s.����D�*4��IY��4��2N�Ѩ��C�}(�8���V�l�F���q��.�����5��pc�������*�� x����A.�5��|�l� An1�.�YW�.�L^O]�n��^	D�O����K�o{�޲�@��_Yk�
@��8�a��S��^��%��6���g�����]�n.�	��V����n|��*�tJՖ����B���9��Vgd�Q��<E`O}_ꩼ����B���o�#-��a �-#jk�Rݽ׾���]����/�dOE�±麸Y�̓�UL����~3}�<��+��,8�՞󥀪�U�mm ��'�ɾ�r��(a�'تSG2$��A���޾�Mv���e������В2��КGKo�K&f���G��q}7��.�F��n^�c&AJ�!�ki�O'�/����������1��^��!0�Z�vyG���"j�f�Ւ>�B2vS����)�v³2%F�b�Ij��N�?�`��_�c��7U�X$����R��w��e����ܷ��٥#vg)��{�Y�s�󇲚��%���|�Ůd)/���El�4��w/��>��2�o㐑�m��|2���V�eȵܤ���������)q�(��,����/@<���[N����Q��n2�WA�$YR9uX�w<�#�'�t�v����e�*h��&�ZxK~��6�;�"W<D}��P�F��cM�N����g8��%�t�M��d(_���+NJu���X�"�K�m0����?�����Z�[Dא��Yq:ɱ},�ŊIf�]�sx%<�#�܋�"�I��6��+�+�2�31e�M���Jr�'��no�d�O7R���2q�ڏ�����8�g��c�X��NC~�!�R��Y�5j�dKA88G|V���@T.lW��A�x����:��ɍ����H�d�w��8Wjo����;��5�z�4����OC$�(�2W�Mu)�&U_噉S�b,��_yy��Ӂ:�T��ͨ͵Ub��[��VQ\�.;+�)����N����]T�c�w>ϟ��n5��B���y�[�/sK�m7韉@��&�SJ<��b�ȡ���!�-a�~��X���9�.�u�g�Z`�n2g:�:o���6���KBx T{f��{4�d�uU��O T��#U�@P2�Y8�y�̷�.�Oa\����.xo��lS�-g�c��:f: ��X6=$_�;l%�Ph`�;�1Hd�@��"z��Ld���Il}d���MJ�@~R��@}���?��c�<������r	p�}��1ka����FSv��*͗������颽��v�{�G�^db᳚�1�x�{�j�T�����M�8�V^2��9��+���SNZ��v��e![{غ�=�C���v��V~����Bσ���nF�Q��:o�BCZg�:�����j<��J�n!�����t���n;;W&Gb�g9���oW꽪|�h����w�)8 ~g��n]C�J�V��]3����U!�|��1�e��q �q�f�7���>�d��w	~�I�1��#�u:�J�;�k���M��p��?1(�� ���$w�e(��h*җs$�΁���~��对3ؑj�kgī�֦q��jD�̴: ��"�D�j$�	���o�)�d���S>���V$�r3?�ﮯ#lT�ѯUȎ���}[�0�P�%1�B�0�d.-I�b�吽�x��}P#[/
<k)��%�����Y�	O�x<{�p�U�W̹~��J�&߸�}K��c~ly(ٌlSSύ��5��N���T"%����o�k`����[��o�IК�A�Ty~ˏ��[�> DR���)O*�8��q�NʹPs7gio�[/�k��e�2�	U�h���n����M��N��8�ϴ�gÌu�^�W���k�\b'@h��y�H��k��ߺ_ ��[k�Q�Џi]�z���I%Q���	���gF�Gُ� E}�Z����14`�h�X�8��]�N�>A�;Gb<�}�.k�a���QO��f�A�Tw���[z`;\JRk�xW�|���F�-�W�ڞ}�h@g(y���T������ލ�`�1C"q!���pCt���2b�}���>�꟎�v��T-y��J����� p�e*O����F�K�����cF�G��C�����V��_��%L����͚����\4�s��"��F�'������gb��Y57�Vt4{�����c]�b��ڱMsJ�C�-�UΒ�������;��OőR�~Bc��qr�WG�����f�
��Y������̇oe�<)�s���(A��2|Bx0�ZO�ޮ�:���K������^�����h0"�:f��cԐQ����yʙ�_A�\XN������%�5�z���'d�lHs��Ҟ%W�O#e��ͨ��]Mgˣ�+^?�Aa�(X�+���;�=��%-N K�xk�y��װ��]���˙ݻ<����b�&��-�����3`�A�8q�iu�
_���<�����U��{Oc�l=R\K����$(�ĩ�/��"M���ܝȭ�>�[�E�"�.Z�8���d��o'�>�ai�HF���o����}��h������S*@B3��k�	l̲Nx���HPe��_�(��6M7;D��Q�@�e��=?H���'[8F��'7�.�O�ַ�R��m 08R��1�y+'�?��cU�F�4�J廑g��g�=Ë%��"b u�/kd~��"*
��j�@i�-��5.��r�{,S�ܜ�y4W�wY�����*=ӫ9�h'�	�[�$���;̹|2��Z�O[�H��6y��s]��j!:��X��E+�s�9^�I�$��^ �P�74�IM�D�M�$Ć�T�=s�E����W���BQ���E�O|a�\�-O���d}G2�<EEH�X:%:r��r�Ț�eQ�,`O�Q��t��쬦�)!��t��X�EA�wB���Y����C���Q���;�z�7w���x���^}�h�ljS�eT����
�����]��|@�e�CD�r�i�Q�dZ��[l��_@�2~
�v��)ZuC���f���:h@Lͣ�۬j,|�gxm T㊄e��!?��ݞ2�6aC�ܘB�j�u�Z!��(b�8���� �d�����z����&��n>�&��)PW��^���{�~[Zq>�C�͉B��X�|����P�b;��{C��	i"j6{��<�7D�D��u�J`+ֆ�o{(�_�H��T�y�i@yF���?dGL�?�g�����&?�v�.���@��I��E�%�n�c�64í��Jc�^��oU�*�c���}Pe�F�ᓧ;vg��\A��(�ɖ�n�p7biX	�Z��	��o�5��0C��'��¼c�3�c\oX1/���/_�w�ހ��3ĭ�pD3}��;�,H6��e���~@���"c$��,#~$-�qfwp�i�Ikv�rAq�-�-�B@��P�^�
ʓ�l�a�?����2D9��a�	`��B۾���JӁ���|��+!��e�_�=��S�@+�PZ$�Q�,�w�t��(�|��`�3g19�gqA+g����D����h�q�#[7�� ���A���Zu��aP�$	��`���	�'�h�,�B���~�k��Vh~m6b��K�k����q����;��%l}�ų�z��0�l����l�#e7O~B9k��5}�ސ��sFɐu��PZA�X�¬���z�%٪*�� �Tۿp��=<A�R�?{u�0(�<���u!�O�ev����S�m.�����%#�̕X���
6�Q{�&�{�����O�x>�R�n~Xq����L4��߄5������H���� ��7B���=ʻ��X��c�{���(O���Ll�'I�rr��ik��$����Q"���_�%Ja�����ڀ-�SKZ��iI5-O���щ!ɝq��r��B`Aſ��3-���P'�w��[]�`a�NGc�B��,*Q)��`�}uY�� _l��ȦAĬ�}�DKe�5�Қq�J�WwU�������S`�}��j\�x��Y���������f
ޏ�Lg���z�N�~}��|"�4W�E���GU�=��|�7/=�o��gl�/Q��?z��%ml�Ĝ=C.5{6[��"<�J˴;>���>���{.���U�'��Š:җFF茊�� �gW�+!����<y���'T�)l|��b��i^`��e����VS����C��X��N��~޻bӈ�^�n���qѪ��:]U��Y$�ܴD{_�Ar��? ���G�V|Nβ���nWO�dܬ�*FK���8�\y�]Ԋ���D�#30�lmpR�ԥ�.(_��40=ƉxS$�23�,����G����)��H+����TM2��� >�HBTvZ%TG������b�݆���\�w�� �ܖ�yd�\e�f��!�6ۋv=�z�������з��E����V��eba�[�w���m�%+�W&��S�v��$�Z�w��%��Qn���(=�\'H�2��N>ҩ��U�_V�2� �m��y��Q!/��I�����eAQ��|�z�Q=#�Ù	9���'�i/�o]�#���'��?KGGNug�ɽ�]�m�LK���f��|n�!����Q#o�BB����/�rsQ_�L�J:��сW��q\�0P�����"~�wD����i�5-����]v�[���7�4ֵz}E+�%`��^C�@�7n��:��
\,�4A�7!X��z� �I�X�ѿ�/�P�E�:ā�{�D�_��Py�����@t�;W�K��q�mOi9���3{2��Wn�.�=��}Z��Ew�OhS�V}:�(��< wܜe�/�Oa�^X��tDF6�Ͼ���'w�?��.o�:B��AU�OF!����Io咼��ŗD�w���M����d7R-T�*TI[Ѡ��ʂ˳���4�rٟ����x#�B�<���������zi+e�T�a��[��q6��@�[W�e�7�
,G������T�X�4�KBgg��,�R+�\=1�	��e{�9����&J����mԛ_��2�5k6��"Y� _��)g-����)BE~�����Z�v�+�?��ů|O�Ӌ�K��O�M=ݖ�K�I��ء�*���-������2u��553ȥI�[��Q�Iǂ3�P޿ߡ�T�$.U�'�8�:fl-���l�2���QE�]����THy��h]I��ޙ㒋�u�te��d�R3�ц�j�"���[�����K�B�����gN�+���:�ʠAlnF�h1�S�$	�� ��m?x�gV+ܚ*��f;��󤕼m!dW�n�P���B�������jH1*�
�[�u�\K�z�G!G�Z�L���k7<����şd�<J`�:W$�S�������"�5�s���ɑ)�#*>g�֙y��r����!X1aHPj�R�Y��,;�蔮eG��!At��!��ϙ^�O/9�.R+#�oik�Bq�S�'�4���`��z �Gs{�k1��O�7�ڤm8�����{yٌ�^���Q}�m�e�����Uo�O�����)%��7�prp����l$I�#�/M�=z^ �%���ĩ��m��)
�=�t5�w(���(�/ǀ�
p��I�\"��LȀ�_�r��[o�!!�v/�m�n�¸�TM����aă�3�-j�CKf�lh)����6�D�Y!���GFĳ�*rE� ��n�ͫ!X�IZ�U��RoXvy�l�.�?����*��Y�wc�
��9Nk���(��/Щk�/���5�at�K{x����K�>���������55NhaS�4K(���T\�4$�h!/t6��S�@s��N}�m��²���������/��ʘ$�iQ�
Cw��y������Z�܃��&�[��0L��X�S~UYX ����#+�i���,;�E��1�[<����O���5��4����N�	�ӊ�։Q�!o�O���K/�J��j�@��F6poH�w��4�9��KT�d�KH	�w[:�w}g�2�\3+K�(B��I+h�Q5j���Ul�M�6�dM�pukT��{�п���"����
-)��
���qͳ!'��rD��/p<B�P'>l��؎�̂@1�X�d�ߨ9��ډ'X�	�()~!	h�@��m"dhZJ� ����C��*���¢����Gޓy��*LՌ��V�QN�!AB���S���KD&��!4kX�������K�nӒ�M�5�b+&�*6��9�j|�R��DCi)!=r��l���$&p�8�!�`H/j7"��i������Y?�;vcI�P,2�j�/�J8}VN����̜
5��c-Iu��Ԫ�c�H!�~m<��S>�\Snq�#��mb	��B~l��K!N����]U�N	�K��f���Sc�0t��8ďڠ����IH�!`+�j�<+Ĉ�'�,5P�-r��őӵ�%�ņ�9YGh���Dj2�g�X���$G~Cpa��Kj���!�]Y��.0z*Q���5q�@�LБ���'��&W��rS�tr�B ������kz�|۾_!-F5�R�`��"}j�����<� i���cE����돡�m2��6P_?.���-.�<�>��Q�ov���ZbJ�	�[��а�Y͊qm>	�ѭ�#�!ڞ�rl��$�	�T��{{��a%��@%�
)R�t��T8+�knJ�^�QV�+/�	=s.���{��\����~,��3Q��g-؃R�ŵ�P/P(c���r�b0����A�B
-9���=���7m�,�@���q**=���x6sKEO���FO��a]'���,�/�>lc�������x�;iT;_���˽�y΃>]��{�xN7���Y(��	���"�ӡ
wSٶ$������ڣYTr����:������;_!6�T|�>��εL���*5~׶�ֶ.�7���k[���"����h� ���ۃ�v�{A�&��z�Ґ]��wY��W��K�+`��_�.���A݆�g����:��$@�Z��)	� 1��qq.�	rE�j��B�a��/FMN㤲���v�p�Yأ?[m	a��g���[��*�> ߫*�@�x�?5�x��1�MTܵⲈXB�`a:Y\ͧѿ@��@�|?r{L�md#��Ps�k\��T�n�|$5��Z��Տ2d���&<�G�|�	��9�r ��Id2���J��H�u8���5)	�?,�pCw�Ώ�]��c�G����̒*A;�J�t����D� �.�O�.,c��	� [I�7MT�t����������G�>�x ����9b_��Yw���Ҩ���U���d��(�� k���Su���v
}zvO��v�p^=�a۴E�T���D��f�п�: ��˽d�=}��i��H����3+��@
Urx���(�<*�]W8�M�(cg1W璐x[_�tM^�V%ʠ����0�(%�`ɛm" �C�o��ݾ����iz������(�o�an�	n�䛥����3ۭ�Z!�� \�R�>t|�K�RÏ��͔7��|ϺR�S�	d����u3�CLIܦ9�a�[`�t�˛hNr(V͜=֍l��Ёn���D��F�R�'),�QNG��7:�,��Ь�{���<��3) �)�K��Xy�H%��E��ޒɔ6"�N/��Is��-��8]�lT��*�p�>�J�qN=SO�9�MN@U�oj�g��]O!�,Y.�s��`TAxPuU�\���d7&0OE��Qsi*t5�֨p.'�N���Y,�1�8��D4A��T�A� �
U����c0����X�V��è'�:��X��h+�sߣ�B-��L_�e�
K��­i�
N�|
�S�n��R��Q�R�s@��(z�֩�`�p$�ƈ�{buj�1�Pa�a )�I�����BKn�evGp]��g� (tHS�����U��{JF,'y@�4����9t0�����*���/�w��;���]�yH?��ܾ�����ٝ�l�k���tk���]0籼,����d0��w�ߔl�]��X���.�ps~�-Z~�(y#��2��b�v���oh?!B��^
u�o����1,������7#��r��L�Z��?S�Y���b�0�����3��fő��{P� �"���f��O}AA&^
-�E�+_3�	2�:��R�g��m�	����Ze���D��S$4��=�xz5w��S5�ǻY�ӻ�(A��߆&����TX+���/|䉘����;�r�q�쟍K��u�c?�N3�ϰ��ҟp���t�c�F��-B6��ܾ�(+͒��QL�+����d<L��{m��l������޴��5?�ӗ
����p��B0��`�f�s�R]:��ߢ?(|}��q�IXs�ۯ�B�����k�v��(�C����oL�T�?u�]�Z�ʖ"�
b���4V���#��a1��:�O��V_x��gi1AjRS�c������/wG��H=G����H��YG���Jx!R�e���a�o���"�� ���5��f�W���TJ�^�|��%����W��+;o�n;�	KsѵhՅC��uϾ������~�r�z�-s_�dwx�	�/q�"��7L��䋶�Q!|�W����+�]�+� �Oc�?-RN-��V�XA1R0�v&�V�>S�ILЙˊ-�<�%饖��&M'�ܛ�w��sw�Q���Nx��NQ�k_�]j�Lu�ԣG}�T�*,Q�C�o8��ޯ �uC�=A��֡3��lo��&2ʓ��iu����bt�*�bGǭnSa�kTK�Ķ�
$�^Bdϰ���q��� �6{Q���.!u"���%����&�S!,�i��8��$��괽���b�r7f{�E��ˏZs%E��aA]Olj{��-���g�,�8~��@l�{La���#����-դ#S�K���敄(<�=�L�#B�(]S�Ul���h�\`'F	�UʤX!�䛛ǊX�Ńwy���إ�X�	�V�i�	�9�ly�4���bC{ A }C5����i���ƒc��(��,����S�T����{M��|�sSo]���)︾N�����Q��"ܢ�V����׆1�f�3���0_	U���~˧?�6�s���tQk4rp�h�&����T���0�B[�������7���J�qf3kf�c�5jw����;�)g��]��b�lYH%QQ�c,xsV�oVN�X�f�i?.��(i;Mv9�|�L�FR��D�c�52�bז�ggX;\�)�TĶ���h�A����.:��_�`g�sU�ՇQV���G
|��`~x�oHy=K}���)�i��Y���P�M���WR+����;�z�-��.�^v����+���fF C�Gס�莊Z8�u,V���U.�T?���υ��Df/��q���)��>�����f�*y}w+Έ%��7���F@i�AU�w���1��i�W v�:��	�vO���jaP�s5>7�.=��*#�b��RW��w<���^� M6���+k��0���e	^�?�*v'��Ev��b}���h�@v�Z�A?>�(x'[	�[(�_�:��s�J^�N��,0E�,�Xb�����:{�e��<�'{�Y�2��z ��W�s<#�q�=�Ch6��� ���W���U�(���(�A3�7m�ĭ\5m��^�,e��Z�Q-	�6\��52�7[��kp��.�<D_o0�5���}"���6��4�q��h�'��<�P.���M�W �d�%���6h�^w��������Y�IkHiz�>��:�5o.,�_����'�4\CVY��W>�9��N�^9k?���FX�JA\lJ�q�>�%fS��xdNb���U���ĺ��+g�I�b?m�T���9qDY���r��>Z�v5\��z1�j�.z��`�U{NF\_��f�l�^X��N>�t�Y�)(ac��TJ\ּN�>-[{,�w���z�6o#���� ��g\��S��(a� s�%f�!�D��`�3J7<�к>.*	�~�3hx��	�[����9�;p�fC�[�>�E�5*�o�$�_������2%��-՚�2��J��~] ���(k�l  ����P��)�%��L:���K�:��&���"m��+�F�M�g� w}UW�)� 38��:����@�R�$>�3af2�}��X�FK��<%;�P��'�Q��$�z�<,S�^v�>٭T+yY�c+�X;��)��r�ڑ���Kջ�:W)�}S�& I�8�<���*ͺ;>�*�](�D��"j�93Bn�w8F���Za"�L?v�e3��sc�|u�S�&����\s�3�?�p&�K �{�%�Dd�˕/`e�<�IF���_[��q�F���K�oJ��E������(~;C{��⡶Ja��{��	�.X/����N���$6����G��G���NU4�M�t��i�a�����l�jm�W6KL�y���	���J�ްa_#	��mM'�������Mq�?xP妄�M��J�f�P��L�J~�.y���h��|6�y�b�>2؈�.��"*��e@0j	�C��"��;#d{�U�CI�;��
��ҁ�"�����(�v����'kړ8ES�:҅�Ԝ�����`���R�Q�[}o�/���������q�}H w�K"�y����Ԋ�,����
aS���ס򇔔����}M��>M�����eZ�FA���.�K��V;b�O�,�Ҳ%��a�.#2�O�$���尙���]����fO
�	܁��TJ�릝��M#�zS�>��`�G��������_N6V+~�}y�5Nǋ��IpS�ܨ���Yu�0�	����^`|�EI`r��/����Z��]yp���/m S��x�G���y@v�r!{@'�5qt$�W&�ߞ��2�9�`6�K��]���ǹwvP?�W_��~SP��ۆ8#P�L��XD��Y��.CYee�o/P������X�+��wv6K��WZ�\��{��X�^��F4�(Q��d�|e���"�Gv�B���m7�R��LO�m�05S�گ-k�?��_�KSy�89Z�V��,7�9�0�&~t�>
gH����\�bG�$`g���}�y�bV�l��	"�[�Č����D��x���}:�x��`hk+b��_���
��� ۲z���w��8�M�
�&�w3J>���<,���Ow�LO,����LU��p�ȡ�v�\zoT{M)5��K�{��W��A���j�ԵX��i�^p��­f�m��DW�x��-2)��}K���a�/�e���[��[����bI�4d�X|Jn1j������s���h�����h��.����0�� ��u�FVja�R�|{����M�E��1?�8�6���8׹�a�����R�I� T��<�2��?�Y�Tg긑(�`�@�m�Χt���	�U1h�Z��.����k�+h%�?9z��!H�骳PC9�[ȹj���ES�t���Z&��#b�����I!����0ǁ	d�3��e����Ê��1�,�pƒ���/��[N���_���� �]l��H�k�4�� ��81�jvs�"�Zam���P�_��Z���7�tJ$�˿b�<.����)- �l��'�&�<(����0F�5��9m
f����9�θ����i�e�?:��޼�Wˬ׽`��mt��ͬ�^�F��I}@hm'�I�w9e�W����Nj�"����r�����A�N�8�tnz��^���lƒwD��qu��6F��9 ;�b#4�2y�z,��/J�+�w�W�j�'�0dZ��%Qʤܩ����u	���g��_L�}w\{����r��>Oa��YB/�	Jwj���1��݁����LX�7���~U�+���VP7�ag�^7�X��Yg.Q˜m<���_ �q��}�a�L�\�1	c;��K��?O�����)o	W���om�ܨLhT`	��K�	��m�M�l���L)�l�]�6���)�D�S����!�*"]|�N$�%��ޗd�K�I2NǇ���%m�b*~h{-�Ʉ�8wMs��|f��? l���r�o����aR���^Bv9w@�xo�OvZY�<���E=Nd_�����gv��$�ˡ���!��4m=B�[A^�α���&޼�ԅ
��{q����g��P|V�/�*����C�A�Zb�n}�z��F ��9ihg�:aM}�eG��p�����+K�MR~L�ä�C�x&G�Wޢ�,;`0���3ֻ���ӄ�����E�W� ��h�>S��~�&�#0ɷ�=��� �i�W�^A���F}��� "��ܱ��q���x5Ƣ��(�AȔX(�S�s�HO��P��	�`-�Ӡ܃D*���$N��T_$b�V�u�M���q�ޓҍN��S�<�S��g�����A����$5��7w�=���`�\�B�o�q�Qn�޽0�b�?��W��R��u�7z�BDoM^�/��@[އ��F��A��wę��K����YtFٍ續����ߡ���wMJ�ʹ+�F�"��)��d<�J�d�d�/J��[;�N]���[c�ͨ���}*�� �<9�Sp�/9�)����e�l�J3����0H	�D����_v���0���3'�4~bܷ��JCa��_�$�\��ĸ̘mE图�����0���	-+Db��nµ�0�P;-�\�0���&���T���e�қk+�; �A���-�Hy��1�#;E]po�>X*��r(@��KFBW��K�/������FB<�R}�J\��p��ά)K�q_�l�l�т�/V[��e":a|�4WT�n�{�JG�;dF8ޓY�D���t��E��K�2��>������,���5��Ϯ Y�����J�h,�cH�e{,-=��Do�9�3����U�Z�JCM4��o��r(��`��e<k�4�&R�	A]<��»%�r��&fZ�o��q���/ɀ�uD2�6v3�{��f`s��b�Z��;r�$p�D��Z���C?@÷񣰕�H����+��E�i{I�_�	~%x�i��ZP]p�'>��P�]їAuV)i���k���3��ENY��O��bkf_;`���/$nb�'�2��"�&���
5vI8���4� �U�E����*���z��sZ�\���w_��wtm!��+ɶY���/1H �O^�׏����ܽ���/)��I�T�C�U	�X=��S����vw�"{� ����F�Z��|?(i����+ڽ.J��[���0$�쀾��Q!�͒����䬪�v	���s)�-��{��Za�w=�F�\�e��_=��h�-��`w�*M�� Ft�-?q�; �)�TO�գ9���;�+l�i��QCYxpy��PQo���(Q3�9+�ʑQbi]!�2H��bϗ����O�)��zn�(Im0�Ĥ��hKE.�8�y���9>�E�y:s~�1��=�U�?ؘ�(G�����%S�M����Z{���Պ��*�F�Y����W�èɽ�c�̤u��Q�&u���Q1fN�D�s�[	�o	�V���ֵ`"G֠RI>|�_v��p�H?1�rB��cL��A�>N?
�����*y���#��/Oo�b�~��ho����,��XI�td(���vt���җ��k�L���sK�����;6w��H����'�%��]�~r��� N�oV� @L�3�T2�����it�ԯ����Q�zu �����ת5 Yj�n�ZA¨Va[�0�=X��bP�o��4}:�C�g�2 v��knu&�6��.���+S8�;kF�����v�h��x��r�t?y&!l0^��A+!�>��5��� ᭍[@��m��.c�7E�,�4U����QN�ȾE���R��dr���q��\�����nq�Z�UI������m�E�NA�2��MК;`�bo���$����R�2�pɭ�\��W_�A��}$���~���O]���������DÏ-׽�R��:К�;���^��(��1W%묇D ɬ�TD�d�:�U��#h��J��t-�{}�?��Nj�󘀼@���NsѸ�>��(T�����y��������n'�s���Bˢ�v%n�o�+�`�ٿ^�>m�^$��zm]f���FE��/�;�J���� I֮�0ې]^���(Y�8pyE�/���A�+���YR�O�j�u����y�4�g��'���*5B>a��cI�����!]�&��p�<+r�>^�[�OWd,��<Y��X��*�t���)�����Y�(��d�8t�+ʎ�����S+�K4�}�ه�� 8t�;�������$/.l7#pº�M�D�TB/+{��Í�̈y��a�+�|�R*q(!sR��/�Ӂ��T6!bn����&�v��bt�nt�U�e̒A����ס�ᬥ�"��L�����H�pY�T9rN�;ߧ�VO��y��iT��<�b����ŷɼ� twD66�(�v��C��L��gȓ��!!M��덠W��Қ�����7��i��`�G9��G6��K��Pg�w������:�x���r�l&�9�U�݇�����w����*�)�v����R�Q��f���Q�>�;����c��$�7���|� ����V1u��8��Ԓ��Y&��B8���u[�B���L�(j|Tq��9�]��;cF3����p�v�7�0�7T�
N��0H�N�/7ԖJ�[�:�����k�ט�m��`���C/�h��y�20?�E$��$�OUf>���G�T�����[��Ƙ3MM��ζ�9�A.p��4D�GvA�rvhe��}k)t�?�aƎ���u����<��\BG�=q�����u�g�޺ؕ��n!}=D�?�d�b	����rp˃ͧ2N�f��8@����Y�iR�@+�b(gp���|��\��*�C-W��Oz�R)e������gwwȳ����{��Ѥ?:���Vjfޒ��X������Pbc�����F�m\+3�	�I�{w�l�#�-K��ۤd�,��r�|�4'���F����w1N`�έs�5ĸ�XV�����ak����x�<�:�G��>�|2iS��o�-��3�o��~��Nʬ:~�l���6��#�{O�&�U7�*�e��$�\�y� �w��o�i�6q�rO@eM���X�d?ս �#��́�ڂګNW���ʑ@`8�j�t���^b�D�XmjA �M�=���{���I&��<M1�h���<I	+�m%6wSWD1�~���D�=Ь�,��]�Py���K������F�H����2Q*�{���vh � ��&,nS��AO%\KF@�2Jw��y��h몶FP "|<�+��`*�0gT�Ɋݏ��n�	+������☐���Ɛ�+5�U�4�fb��=���Cy�2�z{@>�����X��v)�r��O
fF������P��O\M9+�M�R�D=u��A��T!��g�+��њC)X�v��k�n)���l�π��E�p'-N����G���f,uW�H�C:hÏ�Z�7�n�-���I
����fd�"0��nw�vQ�6J�[,��5i��Iv_<��]���!0%&��?�	1#�Cn��{�3zٴ�ؠ�����6(4RF�*�;tu�U��|G�qjȏ�� ,�4|��#γ��ʓ&l�|����9�d5�§�G3Hi(��V���}�s6�7�0
o�O�x�^���c�\��]��^m��۠�������;%fD3���/�"�q���d�0�K~"Rpw3_{�h�q�«�o_"Ѹ���/������T*,�f-�ɨ{h����p&R��N�k�%�t	h��Š*�������X R�PC�˭e�\�+��=�X�C�E��a��xE3r {.�Y?X��?�ٽ�w��9�Rʨ#O�k��y�e>��Љ�N��]f���N�����%��0�#�\���iw�A�m��E��j��~HZiyA�	?}����ej��IWU�^��X�<��0��(�(E�P=M�O~$+V�F\$��"��tBᱽ-�껣)�ς9��K��#���~#h��5ͪ��L�ڝ	��
�;z���f'P`���^��g��������!�5�Y��_�%T0i''6��&��R�8�sRO�ũ\|%��+(t����=���6�W8�˅	:��.��o≚M�F���e�C���nH�&g��)��U"ua�8�2p9�M\3�~G��b��O�HC�W���wK���Zeç���� ��3l������P`���_l��4�F�����]�S)W�����.\�����9D����{��D.��Ꞌ$�+�i��� i�������9!�nm�&@��Plܰ�T�obЀ����N�r���k|�^�|D.�Alq��D�Y� �a�Ĝ�}9�ǿO�n)0��Rc�|!�&����L���^���M�L�rI��q�U�
������������V��T7���q�'۳+}� 5nX6x���|�#zxCI7FO��P�gB��`�U�L����`�w�B0=v9�r��XB*�����v��ײ�'S�Ҍ.�K޹8�Я��T��Qb�I���P�o��L�4�y<�x������
��^���H9�0��B�����Z��0Jd�h2�����F�2���8r��!��Q��G�%�qlAH�%���#�F��]�lie1V{����Vk��s��5j��A>n���z����������x�ͅ����,Z��dܮ�b��;x���0�r� #����ƶ@�R���p�Ȅ7��q����,5zZ���R{4�E�o6�'�(��� Ab�A��zD���X��l���_����I��b��M>gvS�?��	�C�]�݌QpZ���hFA�3���e�&ױ~<�
u�3N\7�hl�2�x�!���PZ�l�lٜ�����c�_�m��������+̅u�M~d��Ӥ���
���8;��3�\�֩�����T�N%�%�*ël>��}��,�>��z\����®]�S��ɺp�[W-��jj[#��|�.Z��Ko�w�S
dY"fy���4X�S��F���(�۠�Zn��\NM����K�\+�r��&��0�a����x��%F�5�=���3/�����6Ok��$�c3h�ݤu���؄��/���뫓�$�:���d���f^>�Nޠ,\�oC�E���)c˃�qn�|���b� m��hW'G%_&�4��D=F���s]!���E[)>�@����{1F�	���3�	y�Zㆰ�y�o�9�|3'�9`�A!��_���Z[i�g��ϝ���_����K�N�"'ТO �K:�#|��Ei�Mn���Z��|�ws�4�:�I�������v ut)ڒ�'�
�(	�J�Ӛ3qj�#�D�6�-��,/"p�
�Z~�'��A�����8��N!�
��]�Zi:���!���Z`n]ԪY�֏�|����"�.��Cs��o�"%��y>pbx~�wJn�	e�k��o��	����w���s�rN��e�d�׌;z���sό��͌Q����ˎ�>�}'0p}��7.�g����s�Ѷ֎4�uXً|8ry�\�}e龎Ȑ��u%0�ֳӵ�(Pm
��Z2$��͘�#����6/k�W�^	���m�<�	���7r@=����˿\�=��?�Ί��Ւ?����}��}�_����&�vAO�*�b��G�F%'h�ډ�z��-gA���.�Z��ݎ������]���R��J�M�!SZ*��dS�8Б���Bi����I(�<x�#��y�T��ЂK$KA����cς�-�CL9 ���C��a�Gm�_d���FlV��_����K�����g5����&�`Si�[���&�R���$˚�A#���,k�+����"�.�WCG0�x���A���	��\{��&�b[J�o�c�s�?B�.G���h���g�Ⴢj���v6���CzD�ǉr<k���9�Һ�)F�[lgz��}�L���8m��r*��o���j�ck)�^^���ܖ;��u�B&yJM��{��7�GkrQ��	�s�x�z��j�z,�聎�n��`����#)"w�fJsE{�Y7��-�u*¾�Df~�/|L���x�:7A���sS�Vu�"�ΐ�Mob�x�R�2~���$�u��g��u���#3.�6��{�Έ^�'�r�&��]��S���$
���_��Ň��]$��[�[9�\�܀4�-nr����.�!٩�a����B��*��L#�؅�	Ă�x(ڈ��Ф-�����H;��E=��P�=x�������j[���ϲ!4�ԓ��\\3��^����iƙ/C�����d*�aL���{�%�(2ׂ6��Ӏ����Gs���>!��}��p�#N&�0f',쿅BÛ�������qX�|�C�����snÑVǫ�	���r@�:�TEhM%?~�����݉F�\O n��a�٠�MmCR4��o�7�Qݰl���fI1��f�#��������ȱlZ���&����LoVxȫ�R��[�xm0.��9h�뎫Fb�$�|Q������E��Z�acdS�)s�l�=�����x؀�j��5���8;픗���6nK|��ɼ2x]��f��+�0lBZvb*�sz,	�fk�_X���{m�|����˅�˟�%�Axo._�I�NP�{(��{�Q�Y"�򈖪N��貤J0:�k�;�V,x����x�*���/�3��
P6Wu�U����Ƕ���T{��Z��)cTI�)� O%�Ś�h\�������ubF�� 豜*x�N0Il
�n'˴uZ��f�U<e=�8V���X�Ƀ����	UJ.H��Ex�G1 �_-(8��`�g�t�И{j���yc��@+�5��|��6g�pq#y�w5n.R�1C�	�\O�M*n�x�6��Y�n�b/� �-2=�mn_��&�57 .˟�`�Dȉ;� =���ЮG�6��E�+��\�r�ˉ�f��|*���q�eP��e���Ɨ�,8�l:�����P+�囵��v��%"	"�bx-��p=�P�ot�����Ab����Y��i��(���(�^?�O%���xVfL�v����y(��X�����ͱ�U]���g&���`F��n�Gu���IB7��	�-��:�3���ս�DԪ�
���D�c��)����$��ԛ}�<y#��?����dģ^Q�L8����}'���i�ś`�L�L.�;�>RAp���M���~�y\����w�m�q�JB�S�U��r|�"ju������#��%��x����Ğ��c�=k���Ú��N@8W�1�]��Z��/�!A�����;����,F�.+(�U�����|�J@/��&D��c��a�ؔS@��$����N��	��ɿ��݂��h9�e���f���O~l����6�͐ʡ
0T�J�qڋ�+���/_�h5�r�G?SIi&���wm�|�9������o�;�ú���_%��''�lƂ���I��C����j,�8��&&�6ϑ�d�ts������]�8�_m'��iИ*�g cA�)�M�=�'����|X=Rn�Iog�~��xD����|���=9ߖS���TQ��[�T�X�}HP�
�'���\�I�-k���C/,��ÊbIV�`���F.��H�F�Pk��c���n?9\QZ����V��n�����ͩ!�������e6�u9sן��1�p��N�4����d��.��n��GRV�`<�H�wy7v��z�o�s��Qj��j��Y��-����e��ڧ���.博r���E�I�OM�9a��2`�ڃ�:>���(Ў�;K��ũ}��O�@�`��^]�-�{��&x�lMh_�29Z��fl��^�x�;^���g�PT7y�,!��{*~�cq_� ���7�7�Ӭq��v=�3�\�L�x���L�$ِ��>;j?��R��XXw[�|��������>�'Yh�FM!6���p6���xfX��Lh�m��	���fK5j6f�i��f��	������8�������13z�Ƅ���� ܭ�h�"����Tx@���w�I�Á��� ��G��Uj'��ь��t�d� F� Φa��ߝ�E��1 P���P�/��Ymo6P��q:��=��NҹcT��3������{���JH�`a%]���`աs��P$��e����9�?S{�/O��7TZI�9�7ϙBt_"&-Y0���"\����R�:�,��r��4�K�#Wg���^����r�COBXN����ؤ[���<�ף�v�)Y���f�zL��u�R���K6�Ntj�����+�\��(��ܼ"R>�Y���\u��le�͍C��1���%Hx0��G��jM��Q����uq3�Xw���>D0�F�mv��+�C�	�i���B^�Y� �-)�E��OV���>7�D��k��Q@�8�����H_6�F�$6��{P^e�{��r�Lq�����B.����r�\�i�nj�Yn��3=V�z�ȇ�]'�|�Y7���wyl=�A7͐|0�_�����0�f	�Z���b0�
�����/,w�׫!�ФԪB��L!1�����]��ow�9@���l8��h��'s��\�[�Uu���1��R�Qj�}Ofx+�4�~9�t�F�GJ�Ǿ�4L��������a�$�UEߪ$����԰�Վ�c֩���̼� ����k��j8ꦥ����\M!ŉRxy�"]Y�C�U!�i�R�6��8������9)ЮCUf��;�6|�uگ��X,%O�A���i��e����I�# ��j]+��l�"(s�U2L����}��ċ���E	����F��>aH��t۝2���VH�4�~v���g�����5/�aBA��L`�J/�e�)�r�5��]�K�z��2<�M4�<ǁ�S�M��i9��]�#��'��=(d9���<y�R��f���{0v�C��Î�-Ck�Ov�A��j#�p~j��3�7��*�����,aL��\Z�j���z�8�q2l�,�L'�����nNh�l�*7�;�j�:�yoRW�e�'C���o�V�3�5��W�Y�Qgi(�2�J���N��#_���9�����`<���ފ�����KAU?�==��>����UtD��`�YQ�WQŪy��~��5�=4R{[���g�J���b(��HxWc���9��9Ŀp���\z*�A��K��&�Y
l�onu�rm+����~�ui���3mP駢p��B���VR!��Y&�Z?�@�&�6��>6|Z�uh�3���p��\Pd�E�ce�^��$���������(T��`�[����3ZRec��ɯRN?���	 ���9ve�V���U�p���}}��a`��ړ�D(�LWG���ּ��c�ju���m1��4�3�^�~���V���d%���?��f��lS%��F��{�I�}_������;90��P�x��]OTX�ǩ��", ��d|U;��ӫ{��6 �S�|��uT�\�-Z���^t_j�}�׍����EO�K��-2����H�@{�fv��d�o�L֙6�tD�^,M���n�&b���S��$�ǋ�*_ W�Q�y>_�E?��u X�V4�o��+��㋈:j-�M%�/cT)�h�����]����v�Cænz1ʟ@���4:H�����G������-p*o��m�m1��Q3�^װ�#�jE@z�_��Lz�s|A�ܮ�O����q
垤���cx�+8�<\_�vsA����i:�\�6�@B�+^����+1)�P×�aQ�\kЅ�p��-��N#9!�I�H ޠ��1~?�H&qS��c�Q���U��/���sZAvcU��ݯ�y�ѩ.�b{�&�
a��� �0|}:m}<�鐖j>OSؓ�<ћ+{J/K(�������7�ӎ(*|���U�ZRp|�ſ;�k�QĈ���`oSn��1���ԫ�v�[��U�a�y�+�`��7��^ԯ���gz[`4������@n�Y�vפ���w�P�FģX�mF]t7��,C+��E����Z�,���yDU��}�#��ŕHN�/ 4G���K���'\��{�1�\o�rm,>����w�7�
��͵���
�-g�n�#����tZ��L8m&0%�&s���S9�RW*y�f��N��bY��O���`�"���5�e�XYe8mV�=�\�8�II��B�~��40�I�X�^��	����~eq�W6�����IS�؊kԲ��>1��.u� *C=i�޺8�~�����<:$�<��Q�_
��<��/`A��r�>��D+S勞����I$u�c*z��?�$tE"���P�j5�;@�ܸ��w��A�ÎDΔ-�5gb�P#�Qi�`�Ѹ�g X���� m�U>�^���o*��yRk(���c0ZT���k1�M4���4qxI���2�/3(,[�ݧ�|�٣�U/�!yU�`]Ea����:H|�U���nda���F��6�n���%�G��H�u��Q�?!�f�����x���J3|��	�D�ZV5��k_o��{O� wf&Yր�}�ʣ~����ٿ�2p��p��,) 7�]vw�nL>$�ck$I�U�w��y��a(�t�啍�96�hم{�jy t����p(�5���<W%Y������}�\�������Ȼ{p�d9m�L�V|�k�Q�	%�!��^������Z��K��P���3v�G�4Ƭ.��5L�Ԇ*!0���ƚQ�>��0']/��Bs{ܬڥh��YSvr8�_����sr��� F�`ZZ��
:h�Q��Æ�j�N���p�`�wv΃�������ߺ)�U�[2��k�Gs�ACZ�2��P$O�=�'��z���$�U����2�(ۑ?�����C����L��3��S�1H�O>C2�~�-��d@MyH-z�" SD�+J��ψT	���V�����M�`O+����n�)7���;kG{6!X)o
�u���,��~��a��ɺSx[P@�}�:�O��8fݦ�?!u9��5*u93w�Ll��y����-��j_��ĨU��E�Lyw�����R�'*�։g��ا� �6��fY�.�P���.�c�`.��M��3Dg}M�g����,��Eʮ}H y"�ZU,a�q>C����ߧ+��ŭ������u�U9�UC)#�_�H�`��Ci�	V�'�Ĝ��1�!��e]�s�����x�~���s	X�.�ɵʝ�>�Ljhʳ$@�:g>א�E��\�t���𛅀�Ks�Q��5��P�*��4��X�N-"T�G}'��OvU^֣��j�z��?�B<�d�B�i��Go�����;��;~������)�m-�s��+L㾯��=���U�G�Fn�b�<�]PŌ[�F���2��y9K��j"H�V�����u'�E~W���oC���i��s1?�o���D���Ve�=�@���)j|'�̋3=���n9�Ib���}���8|��N`a����X/s<���}�r\H�	
��.#�'�nU�W�E�5�$[P���4�x��\��f`9�r�mB韅����"��ٜ�ԔDeȭ���K����
:����3S�6�.����ZV;�m1Ȓ��C�9�74����t�+���;c�+t؎����'r��k��8���m�fN��Z|�p|���S��S���C���m|�����Y�-"�����N]��W����sj�a�%����i(k�5S�to�A�|˔������E������_y�[���;^L^y��,o��%�y��H�xfv� �w�"�0�Ak�Ɵ����i}z�D�B9]�@�/�2���ng���P��O�0�����Ə�G�R���t"�4�#�1�\�޹�`s�W5Ɗ�V��}��GXR�-TX7Nl�!}܆��YE��L(m?�j�F2ѝ<o��B�����;r,7�����pV=&mx�-�c����u�����:MtRվ�rȋ��M{���p��˂HO�[����BJ`�D��u��$U��P�r&�i��xp�/�R����&i�Hf&�'��B�TZ'rl�&����[�+��!��
A���Z6���ս��(Ί���x1|��������(_��L��e%�o��?L�U��7�lޟIH ۲H��A ����yp_�J}k;�ROW���ÎZ�޼#\+�š9�ݷa]P�E`0�(KY�����T�%�9�E�	��D�݈޸���W@�DZX�[��	�Ňr�H'�����`��אi\�a�{F�Ah�`�T���_���n�(�p�gm�*��z� C�v�a	 ?�k\�@�D�N�vc��n�#e
�ke.b�<��>܊�?1u�Ч�;�ϫ�\��L�_��GRY#V&�/+�R���F�]�1�k/2�O���j	�X䆃RYd{�9��2۫M��%Ս��y���V�8�c�k��W����F6�Ɗ|�i�Ẍ�B�����$�����),ڕQ*�u���`��+Y�*�^�vk�B)��y*w�ؽuv�pJ)&���x�M c�05��~D׳��&�I���9ɝ����f�p�-�{g����9�/C� ���v�c5-CÍ��k���,�`]>b.���f�ew�R-����x5�Ƶ]tN��l2�C�[Qg7 ��8n�]B<�2�x�ho�|кHj�+���*�s��A��3�r~��i��m�5� Ȳ��5�nZ�c'�\������h���L �����Ԡ��;a��⮖g7��q����A�!���=[y�X��Ҿ�Gv�0�R�.R%*I�ꢬf�uK�2� �+ܺ�(�%�M��0��{�u�(I����w܁�ۃ�2&���f+��T���>R0����q���Y8�s]W@b�qn��9�$x�?���}��I̄ǝ�%�jH�S�a�f/'�O�BM�9Q`�f��e�&,��`�O�Y(c��f�RCtA/0ͽ��1�p�� hp@ă�K�ş�DLN�9r@J��lL����8�� ���=-+�ƛ�9J�?�K<6�U�.�Q��ƕ)k��qd����� �5HS���v�Fa_���Ḅ�e��-Z����[�(��f"�y-��F��B#夶���LiX00�_v՚�@�w'VG'���W�F*7��o ����N���.���u��^}(8��$�TI�#��4S�Q�*+�=�4��JhI�_������)cO>w*���E�{/X�ˉ��Zn0�\0�E����"
��,�K�bt`����ºh���Lw
�ډ�7��ϨX ��XGM��V�J���8ѳ��>�S��)��Lņ�xK��j糟��҄����ң?}u���tƂ]3�4�*����W��٣���?uVV�/��c�	�[�f�b,���iW�!���Ш��pbH��[�ı�q�
��$Y���+�l�t��EX0:b)�mtŰn��%�)�b��}��8P�܊����ɭR�³N�{~��Cqi�=���q�R�� ��6��H�84�#��dO��+B��T!X#q9[N�A�nb�蘖�����+>6�{/�j�3��~^�� ���:����|��-;}�y@�]�y&*W?��M+����o�/~|�(���|��;f�ˣZ�����F���l2����66����o=�N�/��>E�Dqh��: ~�q�S��E;1�٤���7
���^�����zB6�Tl��_�hF�{� ���t��E~߫��4��a姃L)Za����-�HmC5�$i��д���-��IK�!�,�<i�a�H� �1�'y��(4[=�?���H�CF�^�� ��O,Z��PO$�rќ�J/~���~�U��ǳ,�#=�E�zEoi�Uj�bWmz��H(���EpT �(���VU��F��tir�_�Aq�`��E��.Jп���/�Ã�Pgę�J�g���0,?470���%���mm4RP�u���l^�lvR��6YC���tjw:�w� ��ԁ��������O��������~%�pQ�w�X�H�}ؿ-�Z�u�
`e�bP��<_��B��Hb�p�p���Ա�7�}^o��*\?XC���m:u7a7��"�k�zY��K"Ir�J�r�9�����������L:Κ����T(T_�a0�P��vr�D0��6L���6����r��H�,J��=q��b�N`��#�
�i�u˨��o�%Vۈ��T����n��$}l��3&e|b�ˬe�:u����g�����q�֙k���U��M��L��5�N��Z�Sh0��ʰ���m7��Ǿ��l�em�`$�J�8"��I����+<�%^�F;.�c�
:h�6���=�TS���ڶ�@D��DK{�	&�c���������ۀ�W��Zۺ��`/fu�w�#&��gN��y͈%���&%�r{�0$���{ �G]��2�,��V&S�(�s����=˧l� f�BW��#�*C�1�~,ð�gmJl
�VS��?�iJ�%��V�� ���]�4f(���A�?]$i�
�)�r����w��?��<�&�f����=�'d�S�Jq���W�m�ѳt?]R�=��U�e�#iҜ�q�����i�۟G@�Z�B��{�&�Yy�#\oX�kcD�-tJ����wn$�U��6(��K+��3R��o�)A��qH�{|=��˦�+�U��� ���l�gUFZ�x�$4��O����*7F�89/��걧��s!/�?�Rtx���NE�
T���;
>��4>
����e����NQBJ8qg����[6�|"|�,A���!x	*w�M܏l�[�ڞWv8��9J_�Rަ3F�a5j��;��a��y�	t̘�@|��HͥXP���䍹�Z���)��ѭ��L�a:�B]>d���txQ�v��7��r����e�;���q��1����łr��c�ɀA�OY����]nnOKm܆)������B،BW�#>�zH���V7�bֆ1��	w4����1��`��B�������x.�v�]v������o4yA�Y�3A-|�^��l�g���� Y�_+�,�Ib�+>r��&}G�41f�G|��FL[�O�����4��21�T\D��%"(�d<��E��&:@u�E��J���c�-�$ݥ���߂J�����w4[1�W�y�����Sd7Է���y�޹BLU�O����F���iA�6n����휄�Yѻ���DN��ܤ��ۦ$�c�e��D%��Jl�c��{F�ؚ�/����z�؇��W�
��*p˳1w���X���Cv]p�'��H�V�[�Pu^�xu9=����ǡ+�u?�fk�c�6l}��wVp�DY�1���+�)/Ǵ	r��ͮ��TT:��~�����E�I-xkv��b^�����?�m��7�_�Z�F(dM�Hz��D��.љ`�ߎ8�/�d�_tj��Y���aY�Eّ�2�\}\Щ�,}8VI`���x��YU�xM��;�@;1���8U��q��m��h����{�S,�D�Q��������|7�S�2+�J�!4��)`S8��?½#s�G�Ӝ��Q�f��$�c�����3�?V4,%9��Z�(�v>gqR�(ar�?�c
`��M�p7|�ףҫ���g�[E/j�A����g�k�A��~�L�}�zfr�H�fV��{A������}���_��Ւ�(✔����Y�|͕�Ow9���s_q��탏Z���Л;��Qi[d$*��˴k���P�Rxp��� ��y�*aN���l��03ٺ�k6-��Y�۝�D�jOOi)A8�Ut�������,/���)�c
�K�����_��dU��I��w	�B-mlo���F�\��T�P!�]	r�H�qTe������>�dNN~U�����;�AZ>Q�v���2�5��2i��@���
�([9?����v�DZ)[�`%�A6�����^�Nj�o�+r��d��t��t��]�����Ս3<����W肂�]�	����.����m�P�ʋ���Z�(�b����ڔӚM ڜ�CpH�����Pp`,)��j�Pz�)��i�M����;e�=���}��;���;a�-rÓ�K����qTȚ)�#
+1�^�T6nz@���lO~��oO���Gmro.�6�喗�@�`4IUBq��P��J�n-�P*�p�2�ؗ��j4�u0� �`>̑�Ċ��>�J�<���KfcA �)�U{힃G�hrifO�A����;��?Go�Dαq��R�Cǈ�@����廃'HLBdz�� I�� M` �JLv�iش�&�
�" �7��ʪt>��[���b�}��,,�G}v�]{�)%^�f�i�F�M���t�CA,!l'�p�͉a�ɫ~�P4K���:��2p�P����<%A�U�,��ہ�R}LP��*f�Ƽ���=�����7�k߲��������+~�rŊp&%�l��#�X:��؞s��E��
�q�Uw@|��3�X��7f�M{�Q�����C_n2iI��D~(��s#r�`���'���i�7�a�Ǌk�����_HD��٢�ʿ0|H⢄8��~�j�q��!�*^	���oߐ�Zk6+��%�m�K����$��&w����i7=ك�!T7����/�~T K�D����fLO����(��e4͖��<V1�jz�	ޏ�Bi���W0������"9a}�躶F̒6N%�t;�:��?1Z� �9t�r��X<Ouv���O�{�i�Q΀�!dF{���6��`�B���PUu�H����@s!����{Ds���E-�����h�&%?�k��V��ڼ�o�n`1�V�f`��2��
�Z)�S:nP�d�B&ҷ�>[۸��t�n��ǧ�6^��o0�v�ogfE�.5��c
��C|I�g�/���m�]A�}�`�� ���L��[�&47�����vd0E�jr�P	\�,��5��<��
7Z���ȩŒX����ř��U�J���>�Z�"[�ͯڸm���.OOW�q\�pz�>��O�TµH��Ҽ����x�`�I�ťL�}�����-�E@�X��;�]�B�ȳv%%�mŴp�����/ʉnS�Xo�~1g3�j�*�X0��H�����/`2+p�!�����ad��@9�H�N�7`��e���ï}r+9NY�y��Ԕ�/�6�S��������؊nӠ�X4�VN�I0)�9I�[ ߪ!�ٺRL&zsͺ����)6�û� tN��g���M��v)^��A捂�
I�H�L�[�70?u�ۆ��/{�~}�E�[���8�Z3&/I[��,�����ޥζB؊"����)zn��l�4P����I[S=U�ѷ��c�����"�S��̴(�u"gp+~�lc�غE�Q8�Dtj��g��]��4'>�38�������IH�R:� �vw��hRi�}3����L�R�\��_����u5�i�k|\P2i:��R��}��oO�.�	B��_Jbm�O	�Z<(i�����8���Jf<(9�`��`7��o󒛍�V��D�P.=3��A�-i�R��O��#FKJ���-��_`G�m~�n���ųml�;��/h"_�9�Y�+����W�,�,5��:��1N���Y��D]����k`�T)��x*G����h7e���]�w�Ϻ^�*'-��~Ss�2;}A{e��/����u�x.����5�n�!K�(:he
��z������o�����D��4����p�X`�{)���$ ��CwBJ��oy�������8Bǻ���P�s�R�"�}>�U�1۱�����=�DOʞ�7R~L�t{"�4͢v���$�#�H�x+;p���e?��YP���F�SU@T~)'��M�����3'A��4"�Jg��
K%��G�
?dHS���o���BE\����5e�b�l���=�^���roy/e�X���cgMCcMD����΁�������-
�Mlӛ��UiǿQ��B�#�{����w��"H5��̳ea���f�o�:맗�A������� �'F��s�H-�?����&>`y��a�,6��)Q;%A+�ǂ��֬Ͻ��zK-?�zK�S/��]R��=	J^��v��i�
2EC4�ߵ0�}P8�Y��٧ҕ��8!���_�\ ���!Kg`xQ�� ��]
�}�J�̭B�}�Zh������X��A��2���)���0��y�W������\�0�7�Dz���s��_(�~Hٖqo�Od.���V�����Jh}Ņ����_�ޱ�տ+v}y�Ӽ&5�apR�òfډU�e�}�J>�'�jb����Z{���(V�5����h�'v�Y�aȂ�E��>=��uY�0fj�b��|�������T.�<)�^��^-�\���\%�;�)e�a�C(�yq����T�̛&���2WV��(�0��3d��?*�/A����<�t#�/�1�\������Bǜmsn޲���#J���-R@	x�a�WI|r������x^�Z$�e�$3�L>':�_���G�<1�j�༥z������<��3�e[ۅq��
�7A��"Sa��y��� �p���J��	E-��o.Y)��}�C@Y;�m�BM���ӑM�%��،���gyw���}�a-���B�:���XD��$�Bd����lS�c�5YB�0��=~e���|\q��]���J�wxO��o	*X����[�XB��K7Az�^�A#��H���P	�u�l�����@d�{�Q�$� yUJ�p�)�*>�}60�&ӌ�y��ۗ�Y�hw��rBy�f��3D���#dG��H ��7C����Ԕ�\�����m��?��r5�N�D����c���~x"(#rm�C3偔V�{!������3ٛ�Q�����n>	���"�(�
򚠲����A2.T�A%�`��L��X����o�;���<��9���Z�=Z�)$I�~I�,�&p�аfla��KF�l�_Q.<�L�i��� ����I�'�{ͫ���P���(��x�8_f�g�ɥZ�r^� ����i�_h�K���,����Zƺ?�:��I�@՟��.%n��<�������c��)y/"齂}<���u�b�k|Dp������p�Nm3�a�>�w���1��P�T���Lt��X]85�GI���w�@0�5J�?��Y*,�m`���s��]]�k{����G/Hāۥ��k�T�7,
�Z�H[-���o����T�3Lt�x2Ѽun-�h��g�,���b,r�f��\���9�>G���tn\�5oT���~���*��P��K�<�>p.S�7�&�@J(㰜DE�=__ZW���P⻹����9�DYuO���^�A	:�C���[� ˵��r@V͓�xQ��_\ٳF+D: Q]
S��Y���Rt9f�c\�T�����.��o�g�W��!�]�4��J���z� }c�S�>Hz6dJ�=�͵�"I"�K}3{N�U�r��S,̴[�N�E;�b+�նʺy�9�� ��Kŀ��ts<4&��b�O�B�B�@��l�V5*���?��'�ۋ��
\;��'���}C\V����ڑg��ׄ�c��ᐼ�\��v"`�
�`'2��>�����#�ߤ<�ie��쐶T�)3^F���L��W"�q(�/�nQG�<�
����6"�:�䭰�6���[�&�_�m�?����{P(lS��ʚ�"��u(�|��(,g�ٯ)�nϧ"aC)���M��k�A�=W���ω�̇�ƌ�8$�E������)��%�����L�ޱ�#A�������P�����~PӪ&���x�eO!<�_T�U�|4�=nA<�!�4�,���0���;�/؛�B�Wϕ��Ա��N�U��+����l�U�/5��fQ�K�|�'�`�T(��e��Vt��@fz~=Æ���U!�*ُ������C�����m�V����Y7�~�O�\� ��3�@�B^;��:%���L��M�D�?���~��L_8z��[�+TT�7\�v�1��]9[?��9�7�';'�+R�eC����躤�`w�>���b����/s�Y\>|O�H���F�ϱ�bCtޱ�h��sPد�$�fX�#Md�y���1�W�K����>���YG�΀i+��yx\��%�;�Y�guM�P�c��m����Uׁ�5�L�-u�vSFZ�:��C������Yko�|�H��Z������ /+&���P�@*����F��i��(��𰅩(����a���rs�͋�ǲp����X�j�qF��F芮�D������ܣžf�w�}� 1n�Z����1�Jq�5�I��Ǵh�);>A��.��m�&�DΊ�E��/�O:!q�Fy>n����Y��2�)���bT"��`(�l�8**���q� w�I�0���X6�^���Œ�m�E��>�1��-6mo	@�K�����O�>���b��i��Z�(�y��m��
 JکX�)�L�����iu(~���͕p!JwlO�li3�l�k��O���A�(��L�N5tÆ��z_����w�|C��1�n�&�D��Lu,��7��kR4t��e��s!��*������^����c}�}{����فWv�v?���d����P8)EEV���Y�lr�z�X���wѓ;��mO�P��Nx
 �*���x���0�ǥ�Er���ч
�Tx�!��ڦO^����d>L���ޫ�Z�b�K��+/0|螋�I1��8?���i�d��������$A�� �y�p��o#nl1H3�o-$��G��J��>�{Q��meɱ[�5hΌ�� o?��ҿ�.�T�<TdqSҭ�/*��-_#᯴�횭"��d���nĜ�8��G��VI��-� I�!��4aY	]˗=&����!��fm��8 ��Bb�9� �� V�ؠ�R$�ˬe�ǑRN�^"N��/�·L��8.Q(��k��#�'��Pha�i�&��;��'5� �y���;�9h���8�Ί�`ⓣv�Q���?9[ Ka��.I_��ֶ� ��c`#����r�`Q?�^�oV.�cA&܇�lk��o�!���ۢ��8R�d&�SqTγT�ne�Tɮ��a�͔[ˋ@�x�`|����'�Q���͆�<�N̋�t� E����Vݔ��M坟�S )J/��:<bOci�u'?�x?[l귌�(�y�<u��Rf:����>��~#��B\ǽ�Fd�{k8���`��Z��Ϩ��� ��(�t�L�{G���?���R����cJ�l�,��M@黚���\�
qFi��{���0���kLh!6��D���Ūf��k�@fx�a�IE7(��Y�3�_��^.Y"��&�C����eTy`[6����pP�Jך����$���g
�t�D��'��k�m��W�!*M��}F	���)���'?�T�$�� �[Qͪ�jj�k����V^��J@gK�����f �i����9���/�f��Z�,�v�h���0�s3ra-e�9֟������}gߪ-���Ȕ�D�k.s���V�J����<)��ޛc�S��ú^�xx�ktN%��4-����uLK�}�0�l5����Pu?�7W�n����ЁAe̋���� �)�G;Tw���
 �Q�G��>�w>;��~����Z���%j��b���u%g�Qs��sg�S� �\P����2���P�/=�"��ߓx�ް�������?�[�D��q�J�D��|I���`�O՝�Ǫ'J���n��X	���>q���Õ��Yքu��P��ڪ�!��)U"5M��ZI�n{�<M��T�e��? �$�S�v7������X��[j��t>�K3{��e3�^9uҾ��O����2�p30fSZ��Lʀ��*�`�"rZ2�Yg�'�l��P7�t�g������q������]���R�1q kRR���̔��%�|<��&u�y���-���jM��v�3���5��{��Z���1(�cf����Z�o7��^߻v�c;�P"C��$[�;���8q �!,�ˣ�k�p�X�f`K(7/%�=.�?g�X ^���E�b�=���Zd'e�%�Vm4�F�Kx�G��h3�,r28�ص���bu�#g"qU�����^>@���&"��;6i� S��l8:�9�Kn
ႉ��|E@��N���dR�hc�n
���Tw��.��8��&4.���1g�Ia~��f�<�h}ۧ�'P�|G'��u��mW9�q��Z6F&M	�a���.�U9撗���X�-����w���uSc6,D\����U��WA�@oa��*	U��.$����<�!X���#��TIL�����`"��aPjx����)�ԡ��v��{/�o��{�
��j֮>xz��E�Gܵ�.��.6�}ŰOk��$Z0J.i��.���,��U,��3��YP/y�Z�M|�_\@��&��&��r�?,�b�c����#f[%�sA�6ugӐ��L|�F��� |v}�`�IƑ�{o��릨3^%�E���c���M���[8掺|O�'�e=S��C*]g������'�D�Y���&����v����}�h�REDǾ�O���#�[����j?�|][�g!{�".YĶ9z�Sg2T��9�j!Ԧ/��uC�.xj�[o�h�D��k򄷃H���Z��Ͻ�~�E�����DvD���=D^B+�����QQ���G��q��nط�H� ��Xcv�6������o+�U
�JY8���0������)ņ��s��&h��f���]t5�19>�Q)tkWw��S/o�7�KJd�k�b�6�eֻAXJ�FG<;��l�$�w�0A�m��(�VWm��*~XK�|g�<R���*{*��0)�F�E������!~��	B����.Q�TV9yj�d�����}=�NΦ��l
O�O�)»�u��L�4��xQ�� �/7��^�@��8���V(�l�Cv���(i�k�Y�ڹC�ޓ�Ձ�Ġ���{ȪP��O�J�g��FR_��P��yN�ƀ:`���)��G�M�J�~�D��ys4GeN�/��S��k�/�m���G��DMl�4;�)��AO�$7Bda���P.b��m�
~>�|�N�_TC�s69���"�����&�,�4+�TSO�!.�*]/��R*/��^W�$,����H�'���_��׍�ɨ�n!ݗ���\{k�OU慂-h!3SM!�ѹ�@;a{���83K�,��K��X�C�г.��	o)�P�ǥ̡F�$+�r�>������lg��!9Q�l�.�c�O�������~R��|=>�8�x��C`���4khZ��s��궛E�;	��%�Q��e�m嵚?�׌��0������~���/T�FI�eZKi��*�߳jf�_��w�i>�}d����
g���j��P	u�_�l�x�,�T�	;��l<�h%�q� VWg�s�0�ފ��p;
 �A_�1|��M|x|�+%�\$,��V��H�����Ss�a 2�k�XTQ�A$���^�'׍Pd��<?�t�*>��j�&�s��=�	��y�܉�3�zyv��稽y��s�>���[_��ax~������#��?W�3�������t�T�.Q%�J5=3>?T-���=�s�͐�}c���Ḛ�5��D,ªG`�fYR���un�XF�����w�'H<)LkMp�.�|�6ᴦm厐�����D[���d�V2��.kV���V��Ba�E�\%e�ȌE"���Zm�悕G����+9>)�d�G��EJ����� �V�[���q�T70�)�{��VsL>��y�XxhU��;/�nhd���%�Pw�<���!o��I_��Zy���;�F>K�~��궴w8�Cw}ʺ]�~����
��[�{�т�i�ƷbN��3J����]-�&��Ċ�����8e4\�@�?t�ɂ�`Þl�F@��:	9����)+��*��E�M��q�i ���(Rɍ��(呬�BM�$R��z淭�V�^���/ɱ�U��P���"��K�N(eb�-�6AOcc��{�+�畽w�9��@��Oe�zP?�J`���@��z�=Q(�j�� ��M�$�~�J�ˤ��}��KuʗZ��9>��#%�q�B�����yo^h�e�����{T`�Ta�-��_\����_"��l�פ�[|/����n���s�_��oI�L��e��x`�%p��]Ҋ`�qp�����/��šEO�6��(c��!��2�B�v����9@ÝC&�<}��iꕔ	e���ć+*8�g��c���k����Y�c'ծ���x��!Hv8�`a���ZPJ�*�d��¼_w5�>I���`$K�)��A�&��Q�v��pM���>��,k�lm��ޭ$�F[�{0��$J^�sm��!��8�tzJ �K���zÉ�����ķ�#u�msJ	��9�^��	�Q9@2�쓃�������%E���v��D4=���p�B_�@`�A�ζ�E�~��W�"@R��*E�,/�����I>r���>�yG����`����<&W�t2���1L�\�B�.-󪔍���q�g~A(�[��������;�!t6¤@���ofUs/�bp�L�<����W@y���@�vsx���J��{��λM���|�|�Ϩo%
)�ġ�2������Z���/		���:��јh�`��=e��\P��}�������eVk�Ƶ��k��@m�;ȷqB~��⹶3���dIΝ7�A-%�|���~-�|V�`���c�K�Ӵډ�R4�ƃ4bo�?T�}7���?A;���Tm��b/z%%�����Ap�$u~G��ý����,˘)N �)!)�^�J���|����Y��ߪ6���3�8 ωa����nV �q9����#��e4LQ��C�zR$���Ά�47�$�2�/4����C�t�k
�쩭����Vw
L��5�U�=C^^`ٖ��|�H���){p'B�w!�<r�� �BBݍ�QM�F���	�ylɶ<9�!asI�f)S�/�	���&���oQtx܎)2��>mҏ�ҝ�{����b�ȗ�<g|��y��^u�x�����Y�3��΂���z�$��Z�H�uy��v��.6P�y}��׳"��(��,��(6�9��q�����欖��n���"�g-�% Ū�R2���M��`j�kD�kaf�/w��o�d�������
t�f�@��^��Z�/�����"Mnܒ~ē;��@��q2�s��b��Zg'�-[��cݔ0�Y�'��}.���b����.qj�/u�� ��[�,�T�}���k�B�6�.�ѫ�����/0��}ơP#���b$`�%����[9ΰ`r��R(�т��4�s���Z�����
�q��y�5��h�riR���j��Ҫ�<&�#ͮO�*��X��]TV�穌o�K/;'��t)'8B�ŭuQa��\.G�F8f�����cE�g=�>�N'�&v
L�Jy��O��`W�P�v��m��,˕�-(a�J�薏�c�][���ƣ�!B��Bc
@����&W�&��X9( �x@�p��,��NXFE��0����u@�E�iz(͊����c��8��Vt.Z��P�����кS:�0�I�Si7�pu�1㛐-W�O3��"lU�؁�<�N��I��H%�^����u�-��A��ٗ�K�]�mmp옩�Z�����i�����f>�?v~z�w-��Ǩ1��w;6�ʹt>#�����cww��8��V^���WT�6b��Ye(	�|�8p>��T�_��+B��z�MDBt`��6�����e]��_�U��fS���嬲jI}��1z@ԚԌ��d&����:��%�ӓVj�b��	ì�
�v]�� ���52�O�aA|���b��7�P���1���܂p��gz��e		e�f/���o
|�]V�����P��!�Q��j�JJs"`Ѭk p�����j�����(�]����̲6��$-��w�9zz�_8r^��e��$�i7�䯉h!�"'(�'�-�1D*���.�"������*�0�lDRl��Fϫ�{�`$c�_/Z�S������I�Hp�u~9������e���v �9��6N*�Ԛ)�Ħ+_��$�J�hs�����������UVu9ěD+�h��a��F�T�ۊn%ss'�_
���sD>�
� ;����U�W���W>nO�5��<亀t3�fyqZ^�L.�8�Z>1=U���_�>:Kw���u�,��M��H��kR���%L�N[uT}��ڙ+;�w���-f��Rd�g����DC�m (��p&��Xy��n-g�����L��vO�5�3/mY~g�Y�)��3�a�+���՝�F� z$�fR��h�p�*�;�UB�����S�X�YۨÇ.�j��m7#v�Y*�*��H_�/J����s��)k4k/P ���U�V�ƶQ��a�B�p��~�$�>�����QR�f44'�����=�a|��Bh��J��˒���G���l>���4���E�6�g4?���.T�v���7��y�yKp�)���D��.�����e�����1��? ���t=;oB���1�t*h�#n����3B��o�%Gؑ\mhM J=�ʤ�wD���F�
ᒻj٤`�;F��ց	�d/&�����؞	X!�V ��Ye�f￉\�g��D��~�*�9l���e�q>�zn_� HaΝ�I6=0񆀝%���`/z9.O����
�9��?���� ����04�I���j����]�FL5���#ۢۯ4)-Ӹ6�*l�Q�\:����:�htGj|}Wbc�|�r�/�6ZU�a��ȖԿ�[� �0b�rB6�G
W+@��0R�ή6��꧋�PVo,�<d�C�l�r6G4G̓8�ޮ
��0�A�X;Y`�.��Ϙ��,�1�R���Z9�u�V	*�/�����m��/�r�6��R �������0��Eن����"��s��ߘ�Ī���W_���H�}힕5*�N(��:���@r�cΩ#��1��K`L�	�_+f��>'y�N%j^�Y9����z��T�(4kbt�P���� sn�O��}���O#�'�'�P���JaP���S���$h� �	�WB�/V'u�,^������x��AR�=�ޜ�N�=Lf܄��R�'�/��=nRT�=8Ez����J��51A�׬����<a���=������I��$��Nx�t����M�e�8��fކ*����b�&�*q���ɱ^ʚ�'�8��Я�g�D���P�����>U>WD�ʤ�S����k��"ϻa�t�e$[��4�F����b��f%�4c.�.����G>bt�;Y�/lo��:ӳy��K�����nZ���cxV��ĒR�#I"��^������4*u?�Z����ۏ�� FQ�+��4��!��a=48���I��i��#��ELʹV�}��]�яN�R9�o�^�H����U�ʧ<V��0�/޾�J�X{���q�ēE��h�RRIW��7a��@���"�kqb~$]�3��`�n3R�|��5h�qj����O�'����s�w`�9�!�7����c��(.K�i۠��t�����1"!�W���-�h�2\�6�=�p4���
^!ߍ���L�ڨpA������+��Wֵ��fV�W]ay�����໤Gw朗ڵN�?���H�8�:TN�F��}P����\̼��h��F��$ǢuZ�~󄞫Ó���:�W����� ���'*�r��]O��93���5��qN���- w�m�`�3!��w��O��ǯ��j��~���*	2Ŧ��i�G�Q��_�:��{�*���N� B�(K�)���b�����G�+�jd�(Q_ �Ϛ�3X<fS ���x.꿩��������3�%DI޻=�mt�	; ��&�(��a�)�3�C4\�j׼17�<��E����w]+�'�����b���H�C�o�������P����/1ć)�����/u�i��A���T���+L���5u�]4���)��^��Kh���(�Dk��J2:b�p�9}��T��s�Q��L�K�j)�NģJ��qo;�3H�g�;�����mW�Lƫj�m��|{C1��(Yv
R��&�ˎ��"��6 X��E��u��o�L+_%9F*���������S��E1O���w,u8��Z���1�G5i�LH)����1z��4[f�Gr���7�Ƒ��j�䩐;`�H�9�EΛ��LI���*�V�PݱT�t�/FW��R�ѡ��ŤϛO���2���n3@�n�C�(����D���D���d[u2��x��)=*"��(A���'�הY�r	bc�j��9�-�Ś
�$O��"+�\�C��И����ݜ<��FA)�U�f�D,�3Fz��J`s���y�����'�/Ƀ)Tkd�{l}9Bg)�!_i�
���8���<=.ێK��a<�"T� �p�D�r)5�[�)n�|�F����X~�LE�IQvke_]��3J�Q���B��x"��D	O �f��T��P��V��g��D�� w��_u=2�{J�OsR9v�vIo�ɇzz٘��P���$�Q*|�Q�{]��	3T������I57R�����A�'o4b��}y0}2!�C4G���_���Zc����Ǜ=�n�1�cQ��b�����/(���5��^>8���>�P�rYT���k��� %S̑!w˅�~X��%\h#�aX���Be����(�
)�^Q:,��0���g.�M¶�����+9Q�ѡ���%�܊Rأ��� 7��>j�2',5��~[0<�m�qy�pBTv�i�~pD�~٨\��	p���Y,�:3�Fo�q��$�BsI�IR���������F����Q �,"�f��LZ����Y>)ƀN�p��β�������OJ�&�0��xm�A$d���P�z��u����lp�wJюʴ���~� �t$�W48�6`�2�,�-ru*1]�.r�󧰟m����(���?# Av��U�P}���iV�z�EW\����ҞE�I^TX��˔��������y𣦲�~V�(�[��S�_����?�k��?�(�����ȑW~�Td�����j���C���_/�^a���R�o �B�e@�����������r�����kSα�����E����s��GFh��i$p݈�ۉX���;����4S7�h������mnc������T�#��n�d@^e�b��O�e��V��!p�^�ht^��S�Ǽ>F��fK�J��������1m�����J��%�S�P��q�r��.J��h7D1������mo�Y���Z������{ 0���$c���j�~[u���Paĉ2���u�@���)d��2es=�_V�X5Dr�l�Wm6ؒ���Hr�
ڃo��o�yU���,-9��4��-�Y� pFcsj,�x����4D��Uj��C��Q��jw��ʝ�	j��B^��y+UC�߶3�8��&����r�7��P����m��R�Ҍ�.#k,Z��ϑ����C^"��&]F���[�P�����	�ح�T#��G
�ʕ�ɟ=wpQV.?�����9�X��Rk�@$�lD�jV�L��忏yk����`��/M,TH�Kc��؅I��7hS=~�k���ߝ���l�w�x	L��@�w�
��h^5�bG?n�I�m��Ɯ��>d�e_�^d}8'��� ����M8LH��]%#�.�%���덋���A������)v�+2S��x�x��Lcu*%��"�"uߝxsM��j|,��?J��Ҭ/���jɦbf� ډ�К]O�zT�`0��x�gz������`�w�f�⁎���o��Ig��#�gY|e 2\~�'G"�X�u�^��1C�~E�n;?��Y8( �ß�A�ǳ��7e�ԾH��-3�\>�����$�����M��q�HYS �����k�����νݩpc*7����Ѓ*��+u�{�	U��i:��)�p�gu��P�j��A�]�S�F�n�H�*�g�p���&�e�'��2��1w�_�+b�sy/��B�Fȉ�1r	����l�˯m��pzU&piY;�U�Xj����r�����Ĕ��ắnI��z�x�^$���%5-�^��\~�t5!E��������#����5�a��߉�[���K��GA��Z�]��ū<X[�3���4��_�-�����CO�JQ�Z��ĉ¼����?�D$�	ˬԡ���z2d2К:��l��$��Gd�/8�tJ�`����/��V��F��(.��s�Z��ɵpܕrI,����E~YK�+�{���r��� 3TI������ug�~�G��8�β��h�?U<=%�����6�&/�YDr��A�f�q7�uK!x��g*_�n{���$�!%��.�\���l�@�Ʊ	�B���U�Za���f�\a^�(�3R~��;�-�)�a~e��[MB���D�j��#O����r5E����D�?��o�e�������>9�H�o�Ia:�)\���{����.���{O4�9\���ڈ����H���]���3�<�_���ZU���|V�>�=�G)%*�s| �	�++#E�c��S�tQ:�I�~5���M[UI�Ľٱ�Hb揖���n#@!���t赽���R��L��q%>Ac%Z~P�'Y�k�Tz��f��Z>LBSĶ��x��i�w���q�m�5|4�04#�o��&[���һH�ˢ���m*�;(��e��twzy��_�C�^:�v$5w��s��oz7�x�;z/����u�WٵGw��gE�|��Z��G��C��?o����Z��D�����将��q���	��5>H��W���gU �	M�����0c�'$O��>E�����d��|���ZdR�H�H���\�G������`zt����:V�Q�SYP�DPzNt��"�V���>�;����Y�	��.y<�����W󾚜����d��ڂH��Gb��DC�\�p	�ۭN�6<�֘��r��T�"[��b���9f�#��*���[U[�ހ���AQJ�L;-�)��Ek�!�$�!��:wĮ+OO�Rsm��u�A�� �"QF����$�����.r5
ځBK��g��u�	�/�z�铊�&�1ӓv_��zܙ*�G K��Y*�d�@�[S+����:�S�1A��#\7謣B��]����@�#;����7�q��h�y���\��_J%)qAܛK'�g`�)2��Y1V�TRFХ�>��U)�'���f�AZj��b���$��[i}E	��?Գ~+�)+ɍI�IJW_�RHY�z.���73J+s��M�y�*U����!�x�G&J�x��j�1P��</�csu����b�z�9ٱ��yOH`��g�'��˷��%rϥo�G���W���+�������j�����Ճ��T}�Q2U0��C������޴�������G�Q<�Xߘ�D$������T�r�z�'>��/~ǟY��(j��٣���	�����4�{��E��_+P<"#!��D#bh�#qGz��Ȭ�MT���7?�Nv��2��EG�콎2��,Q�o�ݱ,��y�ΌL	:�#��4���N*dT],p�&k'�M�u�(c��V)� p~D�oy�Ay3ofxN�����ٙ�<p+H�"�ZxeJ�樺�l~��us���J��3���^�=m5�?�v�|�&s�ϫG��@<y���^>����ƃ;���֣���%"����LG����(�v�E(�o__������/W���E?`��`�T�«x�e�#m."\@�1�Jt�������[(�e�JN\w�~n��bd��-�����(��jC{.[3�'�e��47�7 � � T���l8��<�)wn28�o:��gB �z#��}(g���L���QbŤ���K<wQ��o��̳�Q��/#h���{���9�n�n�f�?|�σ�X��� w�z
����J��0��_�uL��)|�s�%^Z��65*d�!��s��휖�S����8��-o"{sM"`7+w���nj/!�kЕ�(d����P�t�T=&T�+�Se*�@خ~o?KVd�p��m�����T�r�2�����L�Qo�\̘}��5��$@�"���%Y��%by�V3��T�E�=��Qp�/�_=���MZ�a; �A���o-�e��o&@!�M��Y��Z�M��!�{E\YW^�p-�&������[+�[1�
���b�R|�>�"=��?��-���d"_72p@��1�O���=�	��-�D��!������@�3N7쌕��;��:�kr=$ҀQvz����T�U�`(s�d�)� (
l���Pw+�	Q�-��k�N}WslM�DWG����ʿ�ϲ9F/�]��NG-��-o�A'⇛,R���f�|�CH�>�Caf���2�̾�p8dy���³���oW"�4��# ��r��hN�i�c��{8�X=p���"����+x�R���aYv�D;T�S��?��o��~�RO6��]Z�m�`A�D����<� {Dr�����#��1���,r�G��쾶��!�(p�l�oh0[�̙��N������755~�1��i@J�#M�a���廞����}���.PG�������o�0/��� �
�Y����U|���"�����@z���#~��r�#2� s����UM��Sp~��
�)��ە�0M�<�ʹ�֢�$����Y��]����5�����`�f��1w�#���%���)v�)>����� 8���u9�y+mu���9��ٳ��]����cX��+iÿ݈�ig6}�m�v;&8.��fɜbK���b+o�H���v�-� /H��Q�w�{��!$G��E9��Z����dD��`s�[��gv��S��Ӓn��}�[R��uIt���;.�mq�����!$�*�8 9C�`�$l����E��b>��*�<ه)pR�G���䣶#�����g$RF�<�L���K�9��f=��C�Ģ���������0���>��� ��A�ftʌ��}woU��,5x510��t��;)��(��ExUř(Z�#|i��0���.&�~g�����VȾ��18�+�a��c"3��B��7�]�O�n�Z�7-�
�tt�n�^J]��(�{F̅|���[�M�V�j���w�ݴ��8�%�xr�$�>z�*S�L���˯���ՠؔ�׏E�-�&3�3d�Qݜ�����y���6A$��l6�.w�ΥX~��O�ќf�<�Ag�E�4�赸4�O�f�e�q!�0��✧���n`Q��D�U{z����0OS�.(�"Q��8Ft~��&���S�'�̖]<�%�x�)V��6�C�Yd�B��$B!"���Qg�F��h&��F�Z�D �7�Ҩx�s��V�2�E��X�oTP$���(:���T1���x��Ry�y��t�ͩ�G9�םb�����G��k�DOp�
����t�GZ/��*��(�L`���(=
���k�������1�UW�z�S�z?M�=D�Ag!���E���Q�I�v����",q��]��W�mk��`?���wwY�ȁ�� Q�H�a��)!�B��Z��/9
n6��L�ho���łX�Τ.[!�5��1����sُ���^�s�R�7\7zU�M%kq���TH������9Y��čF畔d�����U��.��鹿�I5)�.\#B�� �L�V�����(|6����h��$�G3`�҉��Ck�&։�I F2�?~@f-$ɬ?dV�q:�o�7���pa�c֙�ݭq�V����Ŕ�_O���M�]�`�ID�C���Aq��t����3$��*�������m(��Z����C��������*f�����Sمk���w��	+�$S�3,��������ɝ���x�_�C17�`�e3JvD����s���O�:*x�,�_'�<�g�+�N�����p�[oJ���8�1��+C��L���rNɅ��Gl�>%�kJq+�8r,=d��=��I�g�A#^�"_b�9���孹^��,�w�g\��$TNx�F�8Y`�G%��ф���y�'*���tD9�cNGOH�٣ɤk��1�n�u��m�!SiG����v����wT�j
��ȁ�bu��JF|P���B`�'��\_�Y��ذ�z�(�Do��M���Q5��0B�-qd-�I���xb+ز>��3�]��4��~��E�d�i���P3�N a�:.�d��@����?�:^[;�y�$JǴ��|��v7I	�P��F��~+�u0�|�ft�����'f���"\���dk��J�x"l�q���	 n��o��uG���wp�������n=e���zF�ղ����ʝ/�ڤk�k�O���\�/'j9�t�j�Z������kȜr��ٸ��_;(��h�A7�F�5,7'�7�%䁯��կ=5��E?�/^
ݼs���z#�G�fj��5>�ό��;��#Ș��Mf��jq�1�hK[�34׸E��U�}<ɘ�v�4�eZ�˗{TY�?����=���﫤�r�௰�=zr�A�ƺ���`�k6�+@�h������1�K�(/b�=N�<<�E�t��3ޒ��E���:
!`Lt,���Z�Gg�/��FU��U��4����v�v�P��ı�*�r���3�;�rj.����1�R�s𺙾��R��Ņ\�A�]��2�$���S�t�cf��6k_�d�@><�^��S&�b�nϤ2�lT>+�,AT*�h�K-��2�c�hv]�P_sL�1�9��3��g'y�l�O��VH�07�&�YhL�cOsd��F�^����|$$ϨI6[������j�-�_�IQ���'ͤ��(VD9�03���� �A+In��h�WA2�+�C��]�9jK&2@�a(�KJs�x�7�7�e�j�bE+Sh�y��'�A��S���}��mB\� q�{��(�7,�eu�s�_"%>�i�����[|}I.��	�ZZ `����o�[�`����5�h԰�W���.^����]FGM�+l��i�["���;vR� �c�s��ȟ������@��1��y\���R��p���xh9w1oo��Ҁ�B5/��.�Uz^�CJ[Rzff�8������稀�N��Ytȴxaǵ�U�@8����N8%d)&�/<�_%��lkG/Z)V�AQ�'мÐ&�g C���lxp��q�{k������zT��lt˰l��wk�~��"R�L;`��C�+�aK<����.I��9�-��n���ì��҈���ck$׫\p:/�_���i�Dca�EfI��RD~�>��,��@D���^P|��e��g'�2�&M�؇ar���ٽ��E��A;(�an��7��G�z*���̚�u�f?L#v��$&	�z������^~��<�Q@Pm�Y>�7D+�y�Ľ�Nk�K���`Ӄ�a"�ouWP����5V�G=Au���Q���'�u-]@�m�0�#����Yf�h9=6z����k�}�-�9nx[���{2�-r��MN7�\%��O�ͫ�1����L�']��~3��r��u�wA7s�6��ê������⳯�3��:B�-@�`��\rr��ٌ3Gy�n1�ub��
3{nƦ��)�i�����C�5~@�����]�:o�ϲ�%rM�+�F�@��˱�(�ji��yu��}����J+�5�c���!v�V��m�r�*�2�:�D��k6<by�d��$��;�RF*�����d8Z�S�'��G���d�W�����+s�a������7�J�n(�Q�³��X�v-o:��*�	t�I��Rwȃ���ʳ�o�{GT���٥�j�����Ƒ�zj��-(�Ͼ�U����v��.J�[#�S�ߎ^*i�x[�K� ml$ֳmGF��!OU��r!<	,TP��qG�� b;�d��E{�W����x��4:�B\�
0{-�ȍ� KL��kW�0'�/	�
Lw�T����)�1JU��X�$�`oޘ�f-�l�Q�)?�ƘxS=�
�>�|���(���q��|���w{_�r���l$���V�"¥�V{�M�_�F��*<�+>9�n�sV��w5��b�h��^�����%ı�;�N�Vfڼ`H�60��}j����U�O����3�8n�b���N(�g�v���U�(+a�J�x'��r)�ٿi=�*�0�B��;��܅o���#w���<��yO�C�yP���-�����#
���D�E	�3%��i�&������eJ0�}��*��7�����$,o;��:?d��$�s�	����c����/��+-K�Ņ��E�>�����R���܎����Ӡ�z]S#r��������+,^K�S��. �g��k�%�{H�[c��-8R��g+7�%��p�fa�'1�h,З��O>j��2�m$J�$�d�ti��^�Y-��nZ�6�ʹ;ɹ�^,e�oεI���3�p�nKճח����k�˦M�]dP��l�r���X��O;���p�&��zKC⩨�q�������4!����Kq���?�'F��R���׍�v�>���!o�M���ցS =���4��e$����U"I���Ȝ��Ncd�5B��W���q98��v�TA3��B�Rtl
�E��c�zn_3�&W��_�=�b�{�9���V3u�e�'� ����gO�
)�����0Q��MJU<_& �l��u^�m`@[�,C�Q�4�{D_���K����d5�9��u�S׬�0H.kY~��������4�����m���a�`ʹ ���U��q�>��ic�� �.-ºq*��׍#����<��q�#�ΆZ���Y�ExDXK^r߰H'��K(��R�|. mQ��jc�ЩZ�=�*3���+=���T�C[��,QM@��Dj���RyD�~���Q4����z�D��u�vwaLJ������.���1v��}��p�Hΰ�jmUY�j}��z{����
U�������8��:#�c�&H4�a�E�U<��E_0nL�M;��ԋ!,���^\a#�Әusg`���G�id�H��t�a�o��u˕ӣN&P�X\ ��J~�G�)�Jdȡ4.�U*I",p�r1�z�U9b3v�����Ϗ�����Q(
U?��+6
�K�NX�����R��u?F�CC���!it��#�� ��d�����s�2׫h�G���9	���M;�隵&Cp������4���	7d�VFf@e���N����{���e/6`_n��ZƔXt�f�T7�
�. ȇ�5|c�ʼuq3"��:l�����;D���-���qL=�P��b0����R��\s^�����ѕ�ąe�B���O��Y}6L�a�*���$?� ��!�trAz��+���s�����˹r�E���g�хJ�5��gBd��=O�V�2�)G^U�����x������o`�#��o�5�T O����j3���[�
�#�K(�s��z]b/�u;v��.!��B��s��\z��{zR�}9C��ϾW���� �Lx"RS+E�\yaUv���1�fm}&�]|El����m.��k�����R81�:���
|��ޥ-��S3�G�68=�=���jչ��p@�f�I	n��r������ݝĿ�n�>'�SMX�Mr�"c���Wj�Is�G�Y��v��+�>w�y�"i���(�8��f|�H�Wa��,������P�@��H�z �P���M Cc9h���{�Ӵ���5M�
5��a\_��X�/m_�+�.�E?,�H��ڣQ���e�J�
�����s����1�6K�"q*��^J��V�0^�Q��+ʗS�H�)���y�����M(4@x ���x����뽏w�jMHħ^��%��P���s���F��W��h���.ȇUp��Y`��̔P����F��)l�Ȯ7U�,J�]f[i�[�ັ~�(HS�_${ ]`�S���`pg��C%n��gP�N�'GH`�p���u���K�ӄ2��.�{�r 0�2L����~��`�<a�T\Q���g��މ�8�ɩ���6,�h�~wy�+Z�):A��|���u����&��3m�1���
wm�#B~v=�B��D�qrN�f�b/`t�c
#ʱ��F*�(��I87iaV���f ʘ˥TJa���P���o����g��1�'�3��n��V�pH+��]R�*��|4����F2�?��D1�x#FY�T��J�������J���!��[���S����p�4���ذ�@˪T�Վ��P'6�~&%fe�j`XUΚM��j�mZH�4�,d�BB��G.��e�h��\���,�*���i�2OK�Ld-�캜�L��UƋ�en5�?�U������bB�gk� ��n����d��� �e���gK�^��Z!��JU����ϻ'���wZj�Ј�O�[t.=���P�G�%�h��c#\#����[J��m��n!�֝.��f�磵�������DG�J��@�x�\���@��R�o�&��# �Z+����: D�)J�c��%�E���0	?��w�xcƂLE�KW�ߊ����D�z�J��4�(���	��)"lL6.�wCqw�ֲ���R1QO�H���XP%�;���kUZ P%��|ߒG����9�EU���9ͻ6T�1���:/�Z�S��w�^-%uX�L��e_g�v2��_��Sn5�w{ա:m�X�ۆ���g�X\�qB����i�\.��i�C42o�#В�Ihh'NP�^!�9�G[5`��,g74������<�i/Hѩ�?o�{���L�i'}�ij�ԏ֛��2��1nK�QD1x���Xp�Q�۰��C������qcH�b����.rY�ǥ�7@�������:n�O�{���Q9|R���OHv�ʊ��k���"�b��D�π��-UBV��x�_:�
n:3w~�q5tE9�-��3U�rP3_�Bf��$��Evӟ��R;��x��������[��r�;Gњz��	O6���l���D�8��u�4�%�x��8ah�q ˔�k?���EGf����I<3�0ƾqy�E�bä:-�Q�&�҉��������]�~����q�<q�h�ڻ�����!?qI�C�JkB�3Ac�lk�B�yr���	�]'I��Ƌx��J��� �r������iV
��.�U���q�w�D޺k|T	|����75<<�Y�ڽ=��"�W_�c��2Q�:�J�r�M%s�ˆ�,&���/��"�&bU�d}�`|W��������3�p�È�;�q����V%x��o�����w���d�?�fPV	�^��z�O�hg�wi�I✮/�;������jk	���e1��С���2G�Q��t`w�:KџS����_uZ�rz�,Q-c�Q�n�&]P��|�w&+P�:G�̸��-����	c��\�)�=��p !���H7��^�yOƜxu���|4����x{���x�����ߢ��µ�=�i�2�$�jj����S���-�ԓJ �X�V���+ag�v�F,YP�G[��	�OL6��5C �%�_�KqN�tvc�t1����RD�|+����
]'@�.����|����fK�}�5���Q��0�,�<�V�G��[�g"@�m�m�̴��9�u<{°NvN���h{�S�2+��������?��O����`/c@9Is�h ����z�h�o!���h�DP/Wz�$Y�Sr���ċ�'��E.��]�݁ʙ�x��q�M'=�]�J������N¿���w���a�%�:|����j�4�����^�4�7��9"�6�O���*˩��~mo>/1�z�'� �'^��h�+<�+]�j�g��c�⎗���5������ǘP����9��:/E
�^�%!�4y�d��~�J�e��-���ٷMpg�|y乳�W�5��g.H��L��5Űw�hr�������a�"pF�!]�@�X���:� �y�͒q51�~`�`˲3�$���)��i�i짺_��摞e��J��k�TU��t�y��e�oB�:D0����]� �t�l���Ӣ^/*�4�+EzF�¸:�j>=�9�0�i��Ϋ�P�=f��=f�6{5%�&T(sΡpN��>V=����+���U�D�@�u̾IO���降��lJ[/�@:/PӉμ;��bR��M}Y��[����HAq.��5"�ȣ?��q�>f�LpEm�� 7:|rۅ�¥J�b�9>�Ń�����Pɮ޿��*�
�<���Juv,�!���5� &%!��jr�R�1��#Sm�L�����Q���^Nvb|�G 8�פ_�Ag�?"��*�I����>���yjrj�Ww��&��YN�HJQ$��A��^ݵ���Wx��36��51`�/�Q���Y��b6��Ge!��)Tl�D�@�Y��e,S'\r���o�jJ��p#v�d�<�Y9�����xy~YmP�y������>�9�t-�%���S�Qx��
��gN�BP�Nc�;���/�@i��T?y��w�����:�@?K�h 5Qmc��2��H�R�S�p�}�rr���(���kj%�,��!��ɳq}�Ps����`���Q͞�5���8�4�'M26`:Z���*�}J|.
1�J�E63f
�#AI ��V��T�"���ݼsE,�[�������!���=�]U-�S�\}A;b8������4M'x��CK�j�6��@X��*�ޗ�����z꙯���b�,F���Y��=���w�T�<5�(��'#	�NK1jz�ƟxN>�F|�� �v��p�j-�%����D��ޝu�u�H�g�	6c��5*�M��^����8�$7��I+�����-�n���O�x\7_�p)�Z,��cby�<��4�&��nn��M�0�U��Z����8^8��ɇ�!V��&n���	�02���K_G�V��ϥ9m`�2+�n�4R�  ]r����$4�H(|��qL����N������������i7�Xbj�zt������&��KHϠtB�3EEu.�^�ҏ�O��}+F?>��@������D�R>U�k��ʹ�lf*�h؆߀����)�y~���*���+�[��U�¶���է��خ�����͵w!E����X �'4�_��Ǿ�����W�����]�H����m(�)u 	?OE��X�g���e$10���nm�-Ҝ'��d�	���ʶ��yg &�G<��G���2��d��� q3�zC��Qƹ�	5���H?�}V �h~
�4%H���*�'H��&����g��
��v�R�u��n��j�\����8;�7R����%�&2A�	��`	X��1�f���U���MC��䭍+�u�5�<��� ��$���!�I��xR�,ȉ�hc��G�-v3ݭ+�ݣ���va�H�n�-5W�w"���N~k��w�{Ãdv��ŰVz;�?ү\e��X,���I��[�#¹R���ԫ�����n�l��g&����s�׷;��(�%�w�$��*8;�j�S�3d�+g�_��m���D���=I�)�&���W0��V) �6��@f
�[}��g�s��mu�aU!�L�.��,p潜Ŝt^�Fj�{r[%�Oa�Vj�S���7�_EE���6xI� i�~�3�i��V]8;Ev,[.߯P��K[�|��m=�=�"��'R`�v�*"���=8�n��b��?��Tֻ�w��Kb�>���!Vb��V�/��ѕ;�-�娸�X5h�c��s\���%�j�����u��+T#	�,�f�(R�W�YK��ˑ����ӡ�4��:¿U h���m+*���XA��E�E�X�Ip�f䪅A��#���I����f5��D
�l�=נ��)�!x�fh�xe���;�|��l�Y���	�N0K�?�_)��?yUb0:s?l�-S ]�����0L��BMߠ�����Ό%滼x�!|3i����d��0|[��6�����e:f��j6�!!,��4����P����}S{�j8p��X$�R�mn�^�*\U��q���/<�ёx}\���*�U�0�[%jF�̔���\)�O��h/i�(����ڝyO�nH��Gw՗���0���ܙ25uN?�����g�y��SM�j�$�q���CK���e�ဝ�m^{�� �@�9z:�p���n� �����C�a�~\�x��$�O!d��� �Q����*d��ʝ�����+*����_ �����������"����[BO�1�/��f�\��*���k�e�cjy:l��9#�<Y��+)G�+��p
�� |�҇[��í�'\y�xB�<>L]N�������u]n��Ӄ�j��O�e��0ZI���{�"\����m�;��FS�і��u�jf�"����/��\��Q��+�=�S�u�7��8Z��Ҝ�>�d�=7�t^�Q�^;��@�;��(�#IH��ʠDq\���P�� ��W.|r�Ϡ�kCm��P�۝��XզQ��e�"��5�.�D��>�]%[AHԐ&<�kL	{-N	��[(�e�t�abw��9c�Lِ�d`���?B�]�?�%9�;r+���Վʟ�[��|iW��A$[Q�A@8JYx��h�֑fW]���q'��d����t���k�,�_�,�cW޽:�w*>ޖ,��8�b�+�R�=�[�  ��84E��_B7j�DB�����w.d�Etw�
f[(2x�,���y<;XNݨ�K�E�+�g�+�8c�����U��)�]�����P����;���:���(�Um$�Ao�8*�"#�J�.Xt�A�yp��s1%�r�ċ�s���a�rs�\F�]V�0|��5�j��t��n�5�+l��GD�r^5�19�ᧅ�M1�L�f4��qyr�<
���DHZEr�܃�YX��5��.��u3�G5ˠ�p�e�rYA`�v�B+OJ�'��%���\h�T�D�^�y�k��LF�AR�eN��
��V*��Bl}��	�H�^(�y|����>�Qe�m9�8��vh�dy�s�ÓQ7:6N�,|�K��]h<F��fi>LTL��8�_�J2W�i�%�F��<k5$��8=��t�:����8ju�j�ig��u� ��KC 8�p�zL��6��(���S�:\�N��@RBɣd��p\�Ay�n�hUm��K�I������d(�;/r��B��Aq���E�Zת�s#���ڍܲ�*^w���f�w� �~��G�V�Wbߦ;���_� T�p�w�/����ﹾ'�d~�����{��<.�wl�zl�inA,�E��R�v�D�0�n�y;�=����$�Ui����� �m�>����A&��� a��k�&	��e^(̘��ہo׭U�
7��#�^%�w�m�g�͉��<�|@-k?����ӊvK+�٣.ޙ��l+�1d{�&����)�w�ǲ����?1� D��1
��=T�K;���<Zc D;��WIvh��ѳy4�j�3��U �'C146���AV���t ��{QjxvS�/6_؟y���d�w[6�M�B�?����B}nR|W�B�B�S�|HW��o=��0bz�d<��j�Y0{�`����soAf�d^~�1K�=�4�涪;�V�Ў7ۈ�)�;,��ZL����ya��T����"�H`U�#�j�azr�<J����}۟�xF�h�eh��eƏ���ȟm��*�u���O��C�r��vm�\uN�j*�i,�Xv�"\�*Lsb�	�>}��(>��fIBm����b�;�p�eB6�|(�4M��r�!�i���ǼV?��.w>9d�RgWb���$N���*�!�mW�n�0�����OZ<J�f�Wz�	j��*n�C�E���s"���
x%`9X��On���Ch�ȴ�Qv�`��ok,�^��.M	o��Rm}V\ן3�Y��^Ռ3p�;Գ�6͌~��)���%,˷PZB[Zr\���gS}~����N���?V���*ӣH�0��mx��:�÷������:f���B�
�A�:#緗���)�O���C,�|���(�o�H!y���(�!�]�^���_��JʖiQgK���dȴ��u"�����k9����5n�hG�)t������s�6%M��2\�d���To�ؚF[
��(�/�QBZ7a����\\}�����;�[�KxZX�)lU)8���=9#�3;��U�2?m&|�ķ�^JY�q�����Ծ[2o�����7o/7!(^��=&>��h�pL�`IS������A"�yL�s��V"����M�ã%��Ũ���q�<�+�ݶ䴓"U��S
2�{	h &�fx*��� ��ܔ|���@�Nz0��_��:4���� �M�q9���������������_�8�snHǓ?��y��c���3z̓��~n �|�sQP��t�MY6���e�&�&��7�e��f�`�ѐ���5f�=o[M�&6+O����S�B24�,\
~��H��MO�v�y_C�P[����=�����m;,�	C�he&�)�Y�+����;7��do���"2�;K���C�׻~�!�߹���#U2U�&u-~������1�Wۣk�7���V�&"KC�Y$���� d>d���J�/��i��6���zj����5����0O�ʢ2�o���e&u�f,z}U���k�Nf7$�lo8F� ���M�q�V�αr�3?�O3&��M]0j��)����Uϙ���u��!�Q�=D7$����^��|e�}���e r��k5�T�l��a�K{hCV͟t�;��H���`��@�)�)	�C�vUC8�c'��l�'�Ze$���i+�*����9�m=ޜ�(�&���r��k�A�q�`�v�6��ӭ.�����)�V�{O����{G�φr�m�.�b=�:��>|�h��e�&�<�(^s�U8ـ^0��������J�����e�a�,�Q�D��X
�@�m��>'.�Op[ނ66?��~OZv��#����$c���Q_���$Px��tʩ42��ب��iC͒���s�x�� e<��.�U��@V�q�H�X���f"��-�:�����U����9��0vҼ��'Ћ��K>��]16��=�&Lh�f��|>�A���ö���>�9!3��;[u��6�϶��4.�N7e�B�$�|l�����fE���h�[r���Ҵ~��l*;!ڏ�A��O"ߖ�b�Qv��e{�wW����6�.�w�К=@���<K"��Y/�*I�uL��B�b�')a�.�,nuJe���a�qx��h��\k�(���~Veka����!�\�M����-�&���[���m���Ӈ���<�i8v�6�OF�z���&�a{��s��W���ҭҪ�����Ԁ?r���eX9�b�ĘFө]!���lE6�5�I�^	׼�@��OD�)+����>��CkXέ����8����EJ�z�a
l�Q�r�!|�sᴮY�]��i�(���:�/�.��7������\�r!�7k⑆2)�:��^
)��C�T�kS��)��z�{*��}����9K�+�
Vߋ ���B�w��8]���SK�M��p.�/�;��V	��k�6H��VF�*�S�2ML�%o�e���0	�pz�,5?=�R.���tej��� ����� Eh�"Eظ6���/�k���tC.�L�.��G(:��('��ԑ���I_��!WϹb�3��!�-)�UI4'�?/c���<�]�@���Q���R��pA.ݠ��j�x���ũ�s��V��ޜ����^sݭn�� z���`_������T�X$��׫�JH$�H��
1V�S��ntx�@a��|�
ܤ�.QsyC�`"��,�R4�eWA�l�a����<���C"RZ}2|C;�R��R�����\c���{R��Tl$��;S��T�)�$U5V�۝�>#�nU7�L�Q� �"{�l���`��0�;/dwV&k,�"��c|����8�m��ɷ*�8@�I�Լ�΀!�]�{�w�Aj��J"�C0!�RT�Y�����W,��l��|�\�%d�2��G����I�!�r%l��H
�]�P�.
1=�<���=���ե���ޖ�ͯF]M4o�)d]��G�XM���%<���	�>m����nW.������IY�p	�c�L�:�:4�?+���Κ����aZ^�7is#q��%D�	`��M�yui$���w�M� �AA�XW��Igqؽ/h�ؔ�h3D�0�~��5AO�d��5Cy�2����_��W��i5���XV�F��N(y��U �>�I���(����6��7���y\1ƴ#�.�;�Mqȑ>ڰ�����Ǖ`ҁ�
�g�5����������9 t5t�Q��L(�V%���I 9Jd���	E�@������ϟ'b''9l$�=&H�{FZ�&ʔ��VC�P[�m�����}d�J	8m����(F\U(��Y�v^�96�|��@���%qO�QX��C���CRp\�&YX_SҬ
{\���
��n��M�����@�~]�C�!��"��u�YXn����*�q�S�lovT���1�����V!l�B�A�.�8� �Q=��}�8��⎹6 3����(�v9���I�4'\����w�e1�m�B�]�abL���������xAO΁�Oci��k�l\x*�5.5�c�hǼ2�Lz�z����[��Q�E��r��~.�A#������N>��֍��GF���@�)�kg�p���6Q�,�P�522G�/�W�/�ê�_5�*Ǥ��d��$����e���������U�P ��9���ϛ	�Jg��˶y��2(��k�!�T4Έ��?*as��=�+�l�Q����R��E��Ï�Dsq��=�^�O��׏�`�̺tzϻk���܄Wv�B]k��!���/��*^���
�Czb0MƷyS�fm��& �8I|`i���"�r8���P�ʝ�r�Q7z���S�n_O�����pB�Tl�KJ�gip�� �%}���c�Wٚ�	�b_A�W"f�{7|�]�6����XҀA�7�㢇��ejS���a�!�}���w������DO��"�ʦ[p˵�!Ԝ���a���Ω#�7��;��bZ��I\��
�N�#K��V��Ҭ��"4$t�|���e1)�[���ݲ��(��1��Q$"�5ʳ�j+��Es�� �e0��P�j[����{��;Y,�c+��Ls0CU�2Fz�����s����9N�j��}e5���i�j�]��ֆQ,E,ޣ����c��5ܹs��SLӻ%��pNԤA$ ��?��\dR�:��@��C��Q];��@�kk}�c�}z' #X�X}�λ�"��R��q���5��FR�V���|<�����0��}R�
N뛍��5��u�\�#�S��Hގ�!$�!Sa�����@	�'�W遀0r���,ͤ����_�����d�:����%<�ÏW�؊;��svo������Bb�q�~��U�̀,��TR2�p;�ȰYXm�0��M�䪑C!�Ȇ~#6�F��D��"�jV;��O�?q)�	l�J���n0�����J/"��G���3�	�u$�hR������&#�Y�s�_���	؝k�� ��#0��)V�j�4?��=�Mu�FGK=����HN-8W�#��1ŻG��z�����j��Ҡ���}1������uc�q����;<��w�����ޠ����=n�Aj�	�מr�w�|����XK��[@���P�6`�9��1�@�$�0�yr�5��!�ڶ������(b?�͂	��I���G��]F��a���a�����"���S����u3M߳������q�;<q�-�:]nN5�ˤbq�ǂ�h�g��� ����1��
�74���Oz#^�ݷ�m �#P�=��_b�TIp�631E�wغNwg0�{����>�e�%p�v����n����˗kM@3��v�olp��[��&��9��r����]���E�饌�'O��^>	�/YGn�lK�o
����Dޫq��e��-Y5F�УF	����qgp_�G�K��=����!��8�Y�7�`B��8�ϻ�*�=t[�ln5��kJ{�/���T��ohe��	 0�l s�����x>���"߼����*:�<����S	���<�P6�U��%�� ��sgP� Pro+5jl� �[y�V���a�,�s�Rb�*X������6X������=���������;I��Db=+�>���Hd��P,����=�{��}�d���(�y�[����U'ٯ�`'���@�K)�<�3ժ�e�xl�-������s8���2�����7�q�'����Lrw,d/�iʽ�卋�(܊;�̅K�'Oz)����\�U/��C��?����w�����ƛ\��l"�bƱ�_uc\fVч�?����'œ��s��XIO�A������߰�<�s+�C��C[##�m^ׇ'Q�+�M�]Hh��o�;��j'��@}�HàO�J�2����ʈp���k�����.2��aj�w�$� �2�v,����x3\����z� �L#8���#"d`p�9X���>�飘�&�X7T���Ϛi7D�Mӌ��o���Q�Hiuk��F �ό`���Ui{X�Ͻ����]~wZ[��7)��}D�@�6I��	�
�}��ݙ?�7���m]�]�=إ���������?>X��kx�BQ��]�|kKKsj�ꌏ+�f���\.��<ŎQ�(BEӢV5��	��Z�W��4��I��{����	���3("�=�U;q�R�'�ak0NI�T��>%�\�� 7����9'���`~���x�m�����ɓ�֤����X45��R���]
y~K�Ca
�;b�;ҧ��R5d����G��ȥ�&$�R�bP��F(|8BAJ�
���e{�e9|gUA��%�g��S��e  n��b��s�����X@\�N<P�%����w�ϯg����ʣ�n�4ó��.ՠ�(��ĳ����B��S@ʈR���w����6�	1�{���f�\�Z�"F������N6��^�/oV4�l��8�Br�9<��T9�Y7��u)�#� �ѭ���o�Y�;>=�C���K@��7� ��7X�^e��Fʽ������M��������)9�?��M-�3�k�bEϗ�(3���i4�0w.���l�?�z�.�L��y��7!��]���~saw�C����c,~��U ��"���cБ����W��:�S���vx�tpS�� �3ސ_��ؿ�����ə!�aW?�N2�x�m��^C�o�}>k�� *�|�d�����C�=��L���߀O�j&�������`Tk�9oH0ϑ�D"�Ъ�Aӫ�vU�Ϧq`����M������n���t��������� ��H�p�+,F,}QC�UP����f���N*�0�6�t����YZ������l�.[LqgS&0�Ĩ��˃l�,K�͂oeb&R�2�sM\O�ݫF���m~#�G��Wb� ��ҁ��G)>��
dT٥�v�c����������7_A��X���#=8ɛq���]�����.��Ya�a�«���K�yK�hn��*��.��4?��Bj�$5�.��Y�)��a������G�,?Yhѱ�c(�8:g�`��L���2q�X������7v�12��/�o�x=+F�͢V㉡�7��T�-�\�
q����/�Y��~_]��U�r�,�ⲵǷ��H��;�w�k�:�d��R0�1��k�� ��dmA��!4���e��ؾ�~��Y&�&P��?^�y�WդZˇ����Tk(�"�
�Z��?x�=���ש������e�:k���c�hxɛZ�5t��V;�����;@���
��᳀��;�!=��cwB`C��_9��#I6��)C�K�PG�9"E��[�)���| �4g�:��r 3n�R�ޗ�O�tB}k�|�6��~�3m��!6\���-UH�v)��β��cx��|�G������&"R���f7�p�]�Hk�o�YUIP�M�D�����w*0�1�%�c�`�N���[������ҡP����S�#����!!���N�����:��=�PXa)Q���}6��8���"+x`��Ʉr>Mr�^\��L��f$�s�{z~@�.�|P���^��WnK<
  ǐ@Hm�IL����)��������LN�$/�;ckf\u�g()���c�"{�F�a+�@�hټ��ck��@���2"Nr*K����h������R$��w�ɲ��F�/S
du�C�N�&��Ф���Y/`5��������5E�ّ��[	x������X^1���g-(��r32���@��w��6��萈 YH�_�������i�����X���՘w�[Jƻ���0�������y�@)����W��_2J��Ƙ�v��|�ˎ< �T�����Muh2��ԑ䖺�ͥS)��y��A��W:1���3YV߹.�n����Y�������=(L]T$���G'/'��XћB�3�EJ�. ��)��⛌H.�:�OT#������{�ݸǢ,dkv�x{$���=4ZQ{ƃ��EX�ng\����h�R��Q̜�`�]�0vIY���Rf`3�d5	+:;>��́R��l[��R�zX�q�[dgd�v��(JUL7����D�:M��b���>���'��-���W�oP���Bt@A@l�~,1Α�$)���e+�y�������iH"���U���c�n�!�{ySc�ig)G� K����Lb=¼���p��8�l��a���X�{@���59N{H�K�L��m�L9��1��.���}Qv�c����17��o���@�]k�A�K����]#���ͤ�in�'kuy&S���Ăֽ�@�)5/������4A�.ck��������]�.�z�.���$3��]��.�-�DiA{���n��i��.���$b�*�g��<�`��6aڲ(
?��=��]�#���_pH���9�`ij5&�ߴX�}�5�����vAiN��,	�p���a_#���=i���3�OXKxD�@��55�&`�#r3��Q�����zj,��5n5fcE:0hV�z#Aek�E�a�y}MRx]��uj��D�'��3V|��^��~U}�o��z��H��o��ͩ����F%כ���,D����uy�iN���(�[�w���p��#�^�@�N�������~Zf1��:��P߷
[�Mr��]���B�`:xZ�5�t⦊��(��b�P�B���}#Je50�Arn>\gF�����"�C�X���p����MF�RT3�_�#ג+��!�M���Ĳ���f����B�����G��:`���.���#��'\F0���_��&zl�@Q#|^��?K�>��~͖S�r��N��R5q�#�dG�/ݏ�QDn���WH���;n}�G�6�TaMq�'�.���7P�심-O�)s�<Ϩ�)�	{��`C���"�8U�D��BW�*�~؂D���`@�m-�L�>ū6���}�hNW��r�f\�¸��o����	�σAw	���0�b��Հ.�̱
��99��RX�sɏ�rۺ��N
�g�]����
-y���6N�;�~��بm�4I��_�xJ�L¿q�{����7�E=c>��Ѥ9��j����(��V8�vN\����	�=��ȯ��p�`lm+��F�����-�
ud�`��+Z إa����u�ՏH�����Aj;)z�+Ĕ��-�+ճ,(��l}j�V��g|f�Vt�4�d�S �_}�䧍w���Z��ST��&2$<)orq�h(�[���)��	P�ؒ`��Z��e����K9�� �S��ݑ���zp�U{������#�����y�ԇc>-K��U���@���Y/|�Y.��م��ć�0�k��0�B�)`�ӅV����}AU&��E����, ��a�sj:��z���̓o��G��Ї� aj���A�n���/��^��C��/�rk]��-�v_��,�֖�4~?�UZe������s�y�W������5�{�/F����,J[�]���T��H���jK<w��U�P��2Ȼ��H�>U`����+�P�q���f[#��wDn"#��ɺAH�k����������4���ʊ'��챩ظ-��v���ҍZ�ٕ;`,��+G��C�b\�ƮjPi�<���G��蜷�ݞ(�'��N p1O�I�e��D�3�#a�{7{�h��Ln����66K����t[-c����~���x�߸/h�|��р4���oV>����J���Eb�/�	�>�`Y:\Q��k�L��3'U^O ���B��� 7K�,7pRM{֔Y���7�9o����*��Ӹ��eB<mP"�U�KJ&"ޓ��*�:%���Ќ	���B�n�V���M"��i�ݙ-��#� �Ȧ='��ZeI���Q��T��h,5�7���药�.���h/3.!.`?������"�݊�_b�^O[[�/�&�m�� �*.�Z4��?�L���Z@��J���Q]��1�H 8"�+~�G�I$��?q��,�V"q����|h��N3�6�j�8�U������>���7��������r\�1�?��K�ꚭ�0�T��4� $V�ćP���髢�ʏ>�*�o�+��`�v�Wٯ�&�p��	Ի5=�r��h5O��#�c��7�Ƈ� }��x��ߊ�l3�d�hx�G,�5���n:-?5�]z	_�����l娹X���-=��K9��34I�DK�%�����9��?�������DZn���mxPZ^�y��d��[א�xR|	���)!W�HIOR
6@jCx��z���gNu�D&���]H�E*4oka��eKO�*�Ƀ^�m�M��8����!/��'�6�����]�0�6l|�\�r̒D�RG�R/�L�EZ&�.�6�q�YT��̶�$��s��0\dR�g4R�jj�F��8�^�C����8����%�| ��D��������H]��;�	+�>�a"]7����^D�=F�^j@>�W���d�����+ո��i<��]K�Z�?&��fz�(4=�.�l�9�j>  v��F���q�Jw�n��>�N������r%�Z'�"�۞̠a���9M��Qh��������d4EyW��R��~�r���3�:��ܺ4ޖy��d4�2Kk0��l��fK ������3a���m�cm�Y/�pפ�G)%��tg\��Y�θ'��3�4�������eL1kĝY���1�FF([EP5�oX8��fBЗ`��r��j����h�=�dY�qIǅ4?`��~sʙp㣪������v�9~�ٚ��$���;���I�ˇ��"bAt��ï�7��8�� ��$�-���O�cw�%�2�U`�XL �F���E�-B�,���6yώ���o�&���g� �_@�uz �;��5a��:��d��.�te�|��n��C�qW*�F�-8�$\�7>�LNӑ�����`o����U�,h�%���޲+�˂߱��#"���Ʈ $��/?�[�?��+m��8���遛&���Q�ȵk=g^sܖ��dh��SF��zנ�D�oHxe�8��͒���q��ۏ�VfP](�1�7�H��z`<V�#�I�Ql3����p��3Rb�+��e���T���?��f��8I������C(jP8i۵�
4
�E���X�(�Q-����3Wx��*|j}&Mmtn�����VGf�"�lP�Z��SDJ����?Z9���Y��[`��h��$"b��������3���H@��r�*(�'��AR�e�a����G}�j�uk�j�A/�̞��'��@kG/�%c�>&����ZU"T�V���NU�p�� �IS���`���s��,@��1JBf,=�ɤ]T�Jv��:|����X��M���N��ʝ�����u�q6v='��|�p6�`�'����̫j��U�����2P������������%�Y�H;�}��R(ĺԟ�}a�ʂ9h }E̡���C߲R����+����|>z\݂v;��0����	qi�
$'o�^�sl�M�e_9MR�.s�/�*5O<�:	*�NU�����4S� ���`81�K�DS@ N<8�s�#��a�A���&��a83/q��������N��ݳs�ˡs*��}nH�vw���:9�՟��p��zp"#8����o�d�}�=��?oD>�~�����蜠��i2r��,E@�|�?�/H�
�U�;��i<|�9u7ƀ�~`"z�l	+� �v�(F|�➖��w��$Q}'�<3���[I���Tä�s�%�Kw1��KR�7ł��[G��r�Y	[Q���i'�Ej\]��r�3y�SX�3��p�v=)�J����^n�fǡ��6�j%G��Lx*@L���70�$���nߵ�bRN��>���- a1��H�1��
4������4��?�8o�8��Ol�#���p� B\qԀm�𱇽��*y��E�Jr$���C���|:擴�߅�t�Pe����I
�(�c���*�
1��)�K�/�Sv5L��Y����eI,	D���/���&�8���ZB�\��Eh�g N��Ğ̽J+d�U����s��΅�(T�j{޸K@& zb�~ª ��0��d��3C�g�,$W��Gz�?yH�����ʤ����8���Ƚ����y�
��o���"�w��M���Xe�K�l�Ȋ�e��L.3��b���א�tgUP��f�	���b�h~]��$G���u5e��˖�fA��6��
���P�"���� ]Tz������µ ����^��g��������h,�7�`��*�tdm&��>�/���9�zo�[hsJ�r�g����v�k�Di��r�;G�\����gY��M]��9�b0��B��O����{�R^2�P<���V��S� ��k&��}�?����S��M7ܤ�W\���/hQ�,:�����gs��]烥=�����x ���f�I��7k-��]w�b�pZa�Zm�A�	,HW��oj��[�`d���`�8��գ�[�74�s|.������<�@��Cs�I�������t28��4
�����a\��Vu9p��@(��������"@����H=��"{�&6���f�чzH��h�c ��S��$6maq���'`2{��5&#�&G�&��5̸��j��,����s�|��ǣKY��8+�韯�.�))��F������ U;�霩b
���U��3���s�D#�A�G� �������FG[� I=s\rr�f)\Z~I�����\zG�s<������pY��2:9ڦU����z߬����"�����1�05�F��Y+t�3��̊h� Üo@���3�s�0'Gc���U�l��V��yZ>h|���������yU�^�(Ɣ�Ȏr����ߧI�q��r��}�^7�����g� ����Ż8��dήH�w���X 9�o�P�SN�0�4Y^��]U}�s'8��6�c�s,/�d�i�o�J���P=WM8���i��k$��h�&0�J��8���!�#My�9f����ަ/�Y������E�M���R�:��9�7���Ƭf�ò*�t8��xnm-��:��F�}�c��T�]/��e�]����(��#�2vj��$h���e׉�[lLG�Nd7�w��Rx�¾SH�T8���;[�� Lf���FJ0h�����w+�gh��	r�����z���CN�K�Ġ��/�u8�m��Ày�ޖ��������p�����0��w�US�ލ��ں^n�<�
�GM%Õ���C*��D��l��'�Pv�-�
4Ϟ�����pM{-�ix�Λ]��d�<V�a��������2���oj �sWS��FY�DJmH:7�,����.\�%�ǝS�c�G%��_�}n�B#�K�!�N5+t���l �3�4�:2���C��L��Rx҆?�&]f�n����(�6�쵭Tk�E���?�VM/=z2���ڰ����}Ձ�ueb9��D��� e���A�S��'�M؈x����Qo,���Ӈq���s�Lb���0Sw���Ñ�N��XrK �.�
_�ҏ��i�3}!H��<��@�R����j0�WXl�����W�k�Rx*Z�;27l�#C2�U��KB꒜�7��Q���d�J�$=�9�*�%�]ݯF�G�3��_�,�=^�q�um��T8j49
8��?��ql:�t���Xü_r�g��&�帍�*���]��6�� �;� �z0��a�&yx�	�K��/��AܥHI��_��:��<ZoД��qS����lu����Py'�IR�k���Tᓳ\x8�M.�E^:��b�Xߝ��[���!mVI>?'=���\j+^r�ҡ;�������ֻ��ץi]a�4;Q�U�g��Y ���v�Y�\).ܲ���譃�5�#�E	r!�=�	�]$�󠣾q����Jv	DkW�^��rLo�_��� ���j���=�T8�j�
[DO����R�.Iא�ߋ�K����wM�`�W߿w��~1����)�:=f�c��b̘ƈ<�/s�6�L���%�ͨz{� ���՘qӏ՘�J�w:�)GSt�-N[�'C
���S��JFk*ן��]�' �������@y���?;�Ĥ�B\s􉅿�O�]�`���a��8����49��Q	�7�㤇u��e�5�0�ШD)��oK�a�ƛ��7y(�l��{�E���#��URC�OtkQ�K/�փ�)|c�BW�=�)h���q�� �A�cI�H���n��lxw��I/�n_өmòw��Uɠs����D&�ۜ�,x�n���Ц�btз=��`���~]��G�^���y�l��9ٹ�{#����9}^_�WHq��(��t�&�.d��t���>�6�	���q��T^����&l��F)��>�i�{��x��;���lpT�A�Ze�#��ù��	�����C�@������64?�&p����%0�a���B���� -k�i�2ViY|H��~�7���9�I��'�[�+�6��j��)��e��#�����Y6�u�H�&1��hu����\��mR�'���H�h�K�\�}˓y�3k�p4�(�h>�!���+^�s�`�ɖ�猢��2k��m���U���쁨��+B�
7���~��E&14Y喜5a4)�`*�� pP�2�NU
g�v����e����9'����SA���Ti��� �Ūzܙ9o����DZ�[���d���0�����Tţפ�/iK�R���]��������z��2�:; ^�TX	^v~�@���� +<4z�]��b���,�&=�j�[�k������P&�b��rR.���;��E��<�`����ZkWR��NԒ�7`ơm��ٚ*�5`�7�K�5�W� {.r��%���pT����w3O��a������Q�ھ���x���f�I�	��')[,ݛ~	������'j�tĬܧ��E8�}T�M�fרp0 )�]��^� ̹���綀�����`�;����%����.簀q�I��+n��KrE����h�{�Dh}������.\UCm�9�q�	m�ҟ$����"�m����+Y?���
@�g^xћ�|�z�W�%a'N�{G�=��
fҗ�\Ƿ�z�sd/9T���V3FD�<��$嶉�Vr��i3g�m�҈�-� u��h���;'FN�%l��l�CN��1˫��5д�p+�x��� ��V��J�l�!���wAM�q(�
�h���7���w��LP�1gJ(�W�ɹ�)�-���K�W��e0C�6r5�$vD��B����YQ=s:\�V�{��?�kË:�YJ��H��1��C���w������HZ�Wy=D2��f@��U��[.*m��Q��ai��R|�u��H]�_Y-�xb�~�� g�>���KK���d *��VYyǴ$6g� >�|	�������H���eZ�F4�%{�:��ǁႮb5V��O��`~��읅Hr������ȧ�p���A{�
�{x�߫̐��}�&�Z?�� ��b�A'��w��Ǖ��:4��32<N�g$4�^��]��p�M��A�q�>�AoIl[��jBw��6g9�ŋNfХ��>uB����0免�wR���DE�����V!�Zhy�^��;�JU����,Z��n>y�Y�vzN=m#�.� �<��'��i�O� �Aɞ���kXQ�o��3�ۺ��G����BDEڍ�M�W�o���x7M)C�ln��+�ezV�t�S�P,Q	.J��'�A�(d�.�%���4��f�������:CP?�7)�1���l�����u},U>���构˛g�����Ş��2�O�����UX��$�q����Ac�s�Lv"�߅p,̗��C��*��R�J>��f��;،���_����6����5�n`b�3�������w��J>�*.4Z��D�L�E�3�X��6�U-������̸(Wt:c�_����dj}�e}&s�T�WK��ķ�i-�D�nRB'W
*~�+'�p��C��{ׅU�9$:�Җ���ғ|m��Z�����:�D�O'M�
k����-��	 �`,��M7}���*+�c���S�v�:2NN?D�P�+-^Q�ddV7e�`��{.�x^��"�B.���2���f���̴zB <!4^�m��[@��R�w�#�t�]���U.�د�שU�,�e|ۅ����Ԉ|o�XP��$���i_#�`���+zh���ln�Es#{�	��w�S�#��A�%m�<5|�>�cB��0UŃ�R�?��3����T��X�o)*��k5_��L�(���a��X����`nχ�?f�VR
��܁B�#e��ɔ�r���H��E�n�ە�nx&x�����{Tp]�{�|�d��u�W�-��L�:n��c�pL��&ҕ����փ
�i�]�;"r�B����Tl-�]�T0�O���ao�83�S�߾�����Wԑ\�N=�y �����N]z�N�&3�g��z�o
:z�d��n�H$�J�c�D�]<Z5��dܘO0A��<r�Ê:%?�*~8�|�7�����:M���@��3�eD��q0�R��A���͍����k�M��oB\I��3�����g�a9$R��/�5*���o��c�FD����
��༣��%n ]e[BC(��:�5o�kO&����$��^Uiu9�Xsz��
ސ৷CD���j�5�<��P{��X��h����o�{&���=V5��_ʪ�f0�E0t����2����2����� �P�2�R,e	��.�F�釩��~�Y��G�ӟ�A# x���O2b�0x��.��C��᷺���[�7ݧሣ�4'�N��H ���V�jR�$mn����v�̛M3h�!�)i����V,$�w��y�)�+����"��J�7��`�"�tyA�=a�eǗ����GJJ#�i�RG�U��9�̴���3֡���M.�#�m!\�Iɋ�H&Eս�TY��PQ{-�KR|����[Y�x���ݻ�>���ht��}�hXe(Sd���b�:��I����YCP��҂Z�=w�_FƎ�A�xx+��ߺC���"�����T#�f]�BMq�W����Y+����j�\�_YX�`�P�F�	5Y��ӼL�V��)���Qlw�M���
��r8NscD�Nx����!C4�
�& �E�b��8��e��Ɖg��#d�p���iN��$�%<I��t���T��j�b�}�l���jJ�������=�D�ɠ���/&C'4=�0�T�b��#�rh�/�,��h]Z
� ���qÈbdd�q 0�=�(�|��)g������CM���+��Q����|�ɛ�s�D���I̍��s�h�=g05�׼�P)A{��aܓV�R^�܃(��0q;v֑�g�d����X��*})�aj<�>�Hn"i��{�����-.�,�y��MT�/n�m�v��wU�z����V���mEH��s�[k�|P����j��z4}M��Ò �BЮ��]Z�kP2U��gܿ�@�U ��6>M���gx�!c"���&p{/j�c}��Ra=Pp�4�L�cy�7�.>��&�����o9�WO�od�;9������e|KuW�P�0���|�]�dxaИ�F�'9$骬q��n��s��Bg#�
��Jĉܘ������A��1w�5 ����;+o���ֻ0߄F����p��"��皘ß5L�i��#5�j���Q�*���?&�_�����N�-K:D�;�X�[M�:��0�ѪR�%W ���$T��A�C�2�mF����#�fq�*�5�Oą��h
4�����/�a�,2u�`:^` ��ot���ݓ�҈Y[� %�>`�_�>X�XZ;k��q}���0����l̥�����%�1���� 6!H��)�e�tn����#�A:yq���Wޏ�!�:�j�UrH��3]-��V��N��	6W�L��r|b��>��e�T�[n�_��̶hy�q4��ëYyau�F��6D���[�<`�K��6g�|~��ş��7:��l��x˰��i���IQwZL���q03�Y|��t�����%c�XՇ���ˀ��{x=A'N#����m]W.�PϦ�2��G��K� |8X���|��i��Y�f��)|n��a���Y2^
Uณ,5f�z����`�C�^�:.G%K��a��[�7g���L.i#�^|3�r/^ptUL���H���ٿ���O�܂4!j�9:կ��D;��?���MXC���(���_�6�؅�uR1g�l�M�&{g��z*p��r��w|P����c���ʳWtd�<�:n�ds�6% �Pu�y%-3��Sl�8t��L%WX����~�]:�4,(v^�Y
�^�z$9�)&?�!eZ_0���Y��ݓ�,8�d ��o��G��7_�xiy'͓SO�B����y-���e�0Ԗ.��ݷ4Ӯ���>v��}���2�3|N�\�$��"Zy���!�V�ቯ�j�-��Cu6�ܦ�9��� �^]���=��U��e��[��R���rwTo���R��9#bH�S�(wRT����Ti����9����_�
��L�c�C��mH�-t�h������=�2� ?�x�{ϸ^5�� �~=�ר�9w�bp�}�QC$S����n��c��2��(�����VsV����L���f�M�R�
�뻢����7�|�&752'�ѯBe<<i�1&iǲXa�������ǀ�Ih��SR����f3(R��	�ƹL4®3��:�ј��i댚���a�`CH.~�xh'u(@!~�HdY�_n���m��O�l����0��b
��z	��V%�#g��}c���#��1C�q:#�R�K�?u��mR/�E�<@�fŦ�e���t1N-V�-�^�%�J�p�����}	2�g�P�5�c��	��-� ��d�ezo�-j0����'Q��3E�:U��,���\lam�J��R���G���NW�aw}�6����8�-�yp�ǂ�Kq�B��kv�o=�C�}���jz�]�VH�$Vx�� �`I�����5n�J��Z-�������@��z^�Á���2�����Z�U��BRU���B�Q��(q���ȍ�g���-L+��d��5��s�^�r�%��PC����K$wI�H@����ڭ��Ѱ�4)'���;�v�lX�"V����f�̞�;��8�<R��D*��T��;)�p{K��l�%�
���Ơ��v�#�֊q��7�:�"���2[t�z8n���uX_��>�A��	��^�
����=3t~���{����
��z����EU�?r+D��00��� ?��w�%�iC��Z.���b�QS?�З �>��M����dό.`:�5�F6�`���S��ÃI�Ѷ��I�n�]�\����j�F	����.ܵ�� ���r��9�c�I�����q.���a�𑇚�U�hT�R��R�b��s���M1*K6Q�Yk���r�q9����^�ɗ���Y�����`l�x}��y� ��׀�uhtJ0
b׷�a�j]��np	�n͊V�mn�l�4����� ���H3�j�Q��(7��Kom�D ]�4M��nV�ۄ������;�nZ����8~����Qh�\S@��#�����$=��(޿<IOV0����9Glp
��O�鏾w%
��1�P����N�)�ZK��|����z���~��)�<�fM��\�s���]�����:�l��Ng�	�b>�SE���~��|�W"x,t�Ns���&SE b�p�?L5<����`�|�-@�����W@J&o%`d1��)�n沧6ե�f���z.2��w�����ZfK�<�T��#���9����]=����,ų}N��}+1��0��`�P���ް�*�#�؃�s�L
�w_��D�Uœ����m���Ua� `�S.�$�3G>y�=am�p���e�"`k	�^ȼ,*�h�R�Ɛ���oX��̮�M��O�vz���G8�t��R�m�p�e�BK�'����!�-Q%���
���������g�!\��Z���g"�?~sW4] 	Z>;~����遲l�T���;�,�&��n�Ade� ����z>��c6>+��f5��|:�k�o�k�7�u'\�nN.�5��oCOu�P��!���ۑ����D�)
��X�Ã���P+�nQyk�a���d�H�k��lf�Y������h`]�i�/��.����\5�[#qs�4����15�y��*�N\Д`E|P�(���a��2�g'O	M��#y�m����z&��2����-�V����@**��J�? Wϕy�A[O�-Mb_�q�½k��\�e"'�8���c�C3&�:S천[����u�w]=�BS�Ü�͕��E��q�����+$R�"@2�U/yiD�]>Y�'Olh.���k����k�pJx�C��g8���|�2�n�rH�˲e^�<I�)�m�[-�R�"fg;\SIi,'!���@���Ȩ�e�<�:x��-_L��J+��J}#��5y�*FI1�m]���� o���.�E�4>Zg��	�T0b}F��N�1�V�ﯕa)�2}�c[�w�m~؛/��-�{�E�6�Sn��\��9��3�hm�Ҭ���#'[~��Wy&L(Z�LR�=��~�&E��o�5��u��Z�㫤U!��>�&��syM�!�c~w�I�|� ۏ�ߙ�6�0�,����~����Д� >�y�Ԑg���y��i%Q�/�$��t��k�5W�Ly�����{��U�������~s��A�J���Gur������ɹqV�����ݫk��݊{�3��Ԙ18�ck�g7�&��R�^����)A�DEZ�Q�j=��"�ym,�ۢ��]�4ĘYTN'���7۵r��zw�E�H� ����4LW����O8���T��	g���'�"��
���3m3u^?��/k؂sh��RH�.V4ы���׎D
�jt�,�J!��"�y'�F�̺b/4��Ş��@H�3Ҵ��
���:�tL�7gm�x��~S�!\J�`;l�>�߀�RV(y/�Y�2�3�k�P��"�[S��vΆ���)�U-D������r=�q�ﰐ��������â�S�ޞ�U����$)vUckGu֚S�S(}(5��J��z�Մ��}t�5���`��<߳O�lv�+�1@7ł�"V�;�[&�.�҃��t,�#����U:j�f��6�D�e�W��?�%�.�t�����A�a�N?�U�dehW�n�&2�a.:֕�)�6�6��
��{:u�#�F��r�h��R ����ClG�}�J��@�*7�$sYj?b�QP�n�b��X��G�؉qw^ln[(��1=�u��)Jb�nr3h��,N��#L�i~l\�s������T���S8ޑބ����t�]�M�e;^B�O�}�5�gn>-���\3-\���ޝ4ٓ�b>�`I���v���8��vj�pS,ӕH���=�c)���
��QrX���<�>ZV-e��l">��#P�\|��Wx���6|��M�IZ���{�5Y��kϤ�|�Ռ�)N
+���`��/��r|��E�z��04�Z�BC�r��l���Γ��ߣT��i���Q�%ԍ��f���7=��.��6���-U��j��"���'�n������DO�5�9 R��v,��BhAJ�{Z��p�1��������SYH���A�el��)'&?�Ƅq�T�V�q�s��]N��L���\=��!H����y��Wt����#�o8��Bd�ܡF�q=&`��n�a?���"���FTװ 63k��\7<��ԯ�%�:+�ea{��Ah�ND���Veö�kb����p��mZi����^�1$�1K��w�Ncb�+��Q�i@2\3��#86����/���<�hp�(s�$�~���{Npe6�<�)݀4�y?�]���/�_�P���d]�����݈R��1��-ၹ��u��s�g��@E�:R��]*�e*��#V{�
�k���TSUW��}�-2���:{9:�[r�@�ړ�<�ǿC��y�N5b��2F5'���L#�\p[�?6��*t�m�F�f��T@��J�@�f�I#l��eO/iBMfm����������oW��w����^��tb�4E���
J5�m�� 0�	T�I����eB�A��!��s�bDw�f�o�_\�� &�����7�q���'݈� >ea+������I4��y
ac%����ǅ��ōW�x��t�i��zHLn��n3��:� D{�ev��\�I9	ƍ�z��}rq�:u{g݈n��8?)`��T��fg} �G�s��B�:����!��k�(`?�,�|�C�;iܕ����n\1j���'h�p�;Er�c�O8�!��<�٩3,����5�F��T�,���Y�Š/NJ��@��ck#�a�R���U�U�/��yQݗ�9m?�����~M�-�/��&��=�6J|1�&l��9k�F�,�1eo��QTm�����n^��[�2���������9�7A�߹`���t!�-����H�x��oo	�	�������cP����q<�z�{����;�1U܋	^M �]n��⯿*_��+4��t��c�F���Kb>��(y��Yo��əف8��
���3������P�F\�_!M7W����@ڔt�~��z��Z�6[˝�Y���̡��ٶn�J�'|���qS�D�D������C@F��5��V���w���3цN��@���Υ����Q�qnKD#�z��t�H 1���H���A\�l�'b"b*�@'Z!vr�,��������OB����p��
e�4��F�nO1�At����	Y��8������(m�������x�D�1=8w�K\�G�Fx�m�s��F��E#� �"m^�݁��'rgd���~�U���p"Z���a\����T���rr%r�[HZc�`����̹��D �:�`j�`���ݍn��?Kz�e�-v�b�PU���&���vz����1���W�5(hjn��,�Uw1X�\�o���X���,z �{w����M)����/|Mn�?��2:m�w�3Ue���!5s�1����/
�+����;���_�$��B��1������&�a�X�#����n�%!}Ʒ���ʀ]�8$#.�b�\X�ڥ������@f���mQ�\e�o�FϾ�N���N��3��M��?HX�a�ܙ�_�%� �c�{h���/g�S?)�F�($~��
�g�$�3�=Σ:֡@>��y��n�sآs(f���M��MͿ�L1�1\�u��fJ�r�����f]TY�_2���㞰11��A����!%�I�In�k�^{ [��du4ĸ�l�Ũ!?hµb���CS�3Pi7(`�f!%_����Z%�xe��.J���aI}iL�P*_���ⅇ.L���a�Oa�U�#�uڹ}A����1l��q���
�\��1UQ=��9�7��m$ s"_8"`��0L�O���ʷ&�z�]a��I���-��+/� :����ʮ�*�A���3�+W�;�76KWC�o@&j��]9�y �|�$�Yώ����\y��3����h��RUy�<s�ǩ�����7�FcN�>NF7}Z\x�Q�����Є1���
j�Dä�H3ʼ�m��%���ԋ�s�y��{<����x��_��8�d)��?4N�H��_tQH�ڵ�/��7��A5Lq���8�LuǞGksN��Fc���?AUx��P�Sd�	�!t�Vz���o�I�e�>�\k��?�X�(5�XT{��E�2G}seإ*	���q�v�s��7�}��^�BKX2��г�2y�����a�o_� ��s��r�Pdrq�h�Y�d��D�ady�e�S�>�-��F�[x��i�+t�|���4C(w|h��4�����W�s�?����U�i#�)�~?6]QI�݁�XՍ$'L/��Ĳag���a<nt+X��
���Ru��ve�)�䲺��$X���6D��x�o\��7��ψm��_`Ov�9:�(-����@k�s/b�[�?Ҹ�{˼�^پ+	N����^[��_����d;����r���6��o��h�d���Y}����;D���t��Ɲ[���
���9��:��%�D!'��-���	j����s�����q>���/����:D�ܴ-��<�ʆpY�� �W4��v��OD3��
ݨ�ʽU:��V�S�8ɞ������;_5a�g��A�~i�Wr�J#ə�P7TK���Oʬ�5L�Ty�;��ͦB�����B���o��K�E3e�:٘:�"O�1�`��]�oH���P��y,R�PDO��>��=��dJ�m���K>��5#\BH�f��1a����1���w)��tV!\&E@#J��'V6�� #�,��Gp�i�o=9�[t�cNU8[0��ht��Y���EC*�)|@>��2Z�~
�Y/ ��w,cU7��bN0UڮC��U,��>X߆�x���|��g�_�<��X`�G�1�}��চ)sٰ�s���MpV�6 �f���"7������*]� ��;5A�VA��rw��*u,��\�L�a�����c������=Ev+�_x>�G���}�%�Tuy�U � &��'�'���ճld��B��4�;gkt���~����6ZQQ�p��R�!G����<Ő���7�P"���(�p��J�`Nz�$�rf��F�w�S?aoЎT�W�F/Hτ��G�!L���BJ��|�������G<h�?s�&p��$��B9��J�6$�?�}���l��B䕼�{��U��qA�^�YK���pa���=��s�2F�"%� �8�|��w�얩̡b��B��tz����.�鉇p{u������lo��s�T)Df\Ҽm<V9�:�8�&(���@����`u?jK�R-p�x� �sZ꽩�	���{�z7��6b�,C�p���^�xu�h�!����IG�Da�f�Q�$��������L���/�W�N��Ez �sj��`]kF�Iz���Ϛ���(�l��_fJX�r���W�-E|�r�j��d����}FS�Vͦ��i�C��xV�=�
�,�mSC�����f|}I�kxkAN`PҤ�Ɩ����]����]N4,�����i����B�����!�v���Cz�ɠ�{��P�(�G�^�e 
3\��o�Od!�{�7 �$Y���\}g\Ž�������EYX1P�+�Ҥs�퐲k~����(}j�`k�;���|t|���W�ݺ�/Y����H�ŋG<�z��=��o��@�;y�]n�g���ٿ�+Gu�~�  ���fe�Iz�j���D���Tܻ&|ȅA%�yk�}��̐�[3*˃��, ���VΒ3zȅ2��@|�� �p�՘'���F�C���N7�~�皓t����B%��[��[I�ª	���7#P�wSkP����G̨,��	�S�����m=Y�d�J��?� Wr;���
���x��5q���+zqI��MԻ�Ml�(d�ӂ0���tqe����X:�G��NϚ�%zu���A��~!�Լ��I��Z���C��9RO��uy�
�9PiJr����9��h|��!L�w�~4bq��Ƣ�����ӫ��$��N� �V��/����yV�Q�9��;�wv�|<��X�F7F���2E�晟�%�ְSB5w� e# �"!������v����t7J<@��鋿(��B�5<$f���s�&p���|)w�u� �\�U**�7S��a+�7ܿ��=*����krP~�&�{��|(Xq`��6�y�P�y��w����H<�{�:�WF�!���8
�����M��X��N�>j��Ɖ���3���N��Y5ݢ]�](�^��=��;�qF����nj�d4���`?��v�qg���LZab�Jy��:�(�g��EJ6"Q�l �R��
%���;ײm�&�9S��"x| C�Y��gsgBCz�&�j�u%`������>�hg��������~�����W�Z��@b�A�=L_u��_�v��	�ݕTiBi��혪2H�U�y鳩1A~]A�NZ�����;��t�&FiU��rM�V�
WϐT�B�����:�@��֐p?i�G�r�Bv�;# "���m��͡�>|&�C�t�nD�/ I��5���䮻���u+	�m`����#f��3�p����ޝ�&�"��&��&��f:#~ONJ�AcpЮ��\��}r�[�S��h�f���F%�r�4Vy�L�����=a��q�W��[�_S���f_R�W����*HҤ�����;0�+���g���5Y�[�@;ׂ;��1XE�ϱL����+`kT|���u� )��DN��t��紀B��={k�i��G�:�?m����@g��i���[��%�̏���h����[)�a�B'%5q��_3�B�b�SL�0 *����9�rK��6�y%s$����oř��K*9J��C��g3�O��T��]�)�`��G[�m����
��s�m���t�dz�,�;7\���(����-2w�>�df�$Ê��;��k��֞�p�O:9����_��w��x���bM�ݩ���(�Ϲ�PB��d:����R�����;�AC��4�(�����zM��]���3̈́�x�:�ٙP(�χB�����,80��s�jɭD�����������N5�ʵgM�$L,�PT_�?��v�
O�t���<�|�O��u����5$��eB>k�Y;�تםM޽}k���P3F��(�%���1r���G��"Rp�X�DV�x��s�_��:5��o�(��"%ղ����ѧ��'Y���3h��K�sxCK:���[y���^5d�e���)�������;G ��AĊ���4���d݇p��61���B�wu1*맥xy�<�u#�������
kbŝ���lȯ��G��2{`O�#)y/�S��
�HmH.���w��i]M����-�)�<,���ĳ����U��q*]|S�:����
�oV�}]�W�ܟA�x.���£�x2�m��j�~�嶂�=�����<鑇��.<�3_�k/bW������5�66���7v?���4Wا�͞�p��]:OM{�����Oj���(����������3���E����=�;���ܚ �lyh^N~�z��`v�(�C����b�f��܌5N���S�����I�Q��� ��
C08�[wqU�6�OAE릢����|�{w�5B.���1��ޘ��֯U���2�Lv��]�'q�]&H�T��a7��k�u6?�#�p}����	�!��]�u�9f�>O��i����Ud��*�(�M��.�$VQ.D#�ݎmZ�	i4/p��y���=�V�g�j���}e�QRQ����2~9��;�k�����D��3���F����:�r��rV^�О�@`f
6�^ۡ�z�\�����%^�fKa�3=�֌~���a�����I|���U4�Lc[Ry�ݨ��+�c���:?i���Dوn��8Xr�:��Moe�?18��n�fsO�YKRW����J��W������l�N��^ֈMvݻT�G�Ȟ6%"S��Z�.�JǮ�h�2����WK�V����B�������R�O�]/=�q��t��<w��N�@�Jӏ!�Y>�(p�D��+�:�PCJ�ÐU��>��t�=���g�F��{�"��+�����"2b�h\��J�/���(Q��:�h��&p�>�����3%��{�SZØ<�?�ǡXP[8:/���tSb7+��n�����"���J)��;U�2[.����0���햏zpi��4�@�����_����ڈ���?<��N��{1���K�_B�̺f�����-;u�42��D���Qڅ�T���v�wt���;?z}^0W���9��r���)~�|cᚊ�]���Vz��H0^�L%h�c��3 \,-G��E'�AvJ:�U9C� c2�󌊴�Ly�샷=M��Ea|�I����6VM=$�j1%>��?��LE������'w�2!�h�#<��۠���G�$<:لE���Ԗ�[dAO���J��Ն���(�
�[��C����P�y�������Y��V��A��W�f`��0+��0��Yl����.ro��v�{֐2���`XI�U.��L�T�����dnhr@����G�ϼ/xҴq&�
҂��!,`�E�u&�m^9[/��k���;�!��3�J���`x=FJC�����M^��D��v�E��"�_˭��f���lW�0�����������|~����Km���!\_ۣtR>�J�N[��Ѳg�"� dʣI�^x ]I��"�iF]���F�k�c�
��8̕I���Q�N����z���vڔ�-/��L#�ki�7�4�E�u}�d#ֳq�C(h�{h�X+���_O���E�P��Ȯ�DMdj	F6��j�uz���s��k)F�ф���R�]�F�p�"b.|0@T�(�U��E����L�M�;��O`�6X%�h�U�@�;ɫ���*��&~�{{�%p=j�����g����	��؇�ڬ��lg�3�|�,�z����V:a���˔�Q*���%>�?
�&�Gw&3O@A���~��^�"
Opeo��tT�Nx{\�����}g��((H���ׅ��%W�a�F�?�t`���+���QD��Z���w]n��2E���G�n8&�n��� �W���^n.�z�����-�.�Eb�k��D�
rzq�R[JeY!�Ej�\7�}덋��z��.\�"�cS8�K�LY�>�����,.��w��%n�<h�H7���0-.����Dw�Β�54'�R�����`xb#��=h����ĥ���vʩ�7^����=�3=���s���䤇�9�p��^ �����'i��`8$Z� ڻM���=�<��7O�粏A~�L�*q�j���c�O �N�bYI�u��ԝG��/��a�~m�����'���uJ�wr��&Rt�@�+��B�i��c%�s�g�6`�ʌG��<V{�:�ǵ�~YȢl�sq�^�6����FX�4G�_$�E��ݷiѯٞ�F���D��ӻe%
L�����X�4��f���r���W#[�֪�/���$�r�����V9�'�Uf!Ȗ���d +���Me6�q��=]��|vW��h9˄.�� Q�}�����	��N���`���؋t��ؐ(ĺi�>�bb
�_�]�I�x�����I���D�,+P3�%m��Jz�2C�ա|DTb��h� ��8���0�:��n��@d�?�Tu%¸Arcu�1#ό{�=ݟI�Rk�h�>5�5�oR 8�GN�o����!���!}[uH�7��(DGy��X�u��m��%R�$��l*>�`����d�0iTx�G?S��s;"n���˟�������g���An�$*u�d�g\[��#��	�۔Bނ[E��%y[���i��&���La%?�R�Pq��#6���]{�g�ru|��9�<>LBw���'��%j�Xc�f�[�wp�&d�Sf{��0�j4+�\��__�ۣ����ʩH�Lن<�I����c`���Q�B�Ă<���T2p��������n����W��˽��tL��l�� �=���G��"�X��� ߎ���+x�Z�����n�����+B�f[�U�t�zmW��V�q�1ӽ�@��p�,��4[��_�	btAm0�ч�'�C8�>*<OWP�t�s־ߛ�ltA(�(a���,녟��3!��姷,	��+Ӱ�����JQ�|绽����$o[}�){B3	*By'�֝8�+�A�>Ȯp�&��F�wj�PG�@l�8�������:�\�����%�t�,Re�HE�Q ���f��V����j��C����'R�&MC��%� ��HX���e	� ��꿥�+�i��b�]k(�Q�E�1�0�z�P��}l����T68]雦����tGYQ0�b@���w���W|�J+#L�	�F�r(�����g����ްS%�(�K���;c�*'�U�-il�{�0����,�� �<K�O9.|�� ��hX���4RxЌR@���=�C�z�YN0��{illi.������m"s(6i��n �R^5�@}$g�_c�ϓ�~'ɼS�6ىRl�2T��T��#�?Ɏ��3��¨h��J ;��/B�Ӵ�	��k�)�`6L���}�o�5?�+7ĤRf7�Q�j��Dr6����*��9?�c�; �vN�
��e��Q���1�3�W$�5j�k��܃�C§�݅��bdhB�Pķ�Z`!��#�^���0��s�{ �>���U5�`%��SS�^�OD��5#���2�����'٧����������eiŹ�~)���K.�[�x�>��Z_���٨1��mu�eN ^!l�O�`c]�Ab79֊C| �=ge{C�v�Țp�woGr�+�/�R$d����Lq�_�����\yLi�r�m��=/��慕�<�9y���	��GO��h �wg�t@�mK$�ř�Jo_��.M3�sZ�������q#X��+�ꉷ.�<ZN� ��
͝ak>���I]���x }Z��q�Nv����I�)��ig0��l5��$Yf�~�꼖�W�Q��ӹ�E��_�a�'5�|���q@��Vd�3:��R�H����\Z����d��y��!�do�J��N�.>���o[y��!���(� ڦ����=�f�E�I���x���X�`�Πy����ٜ�>bJ(>V�x�������>���ꄖ}[Kw_}��g�dX=!�|xڢ6��s��-�ˋ�tx�Q�i����MM$�P�HĨ�S���C�!��8߂9��)�2ͩ���Ѱ\���g��Fr�����5	_�{`7'���������h14��t���'�en2���%����J��֪��t�<��;�;��j\�b �nh#�n0���n����z̳hj��b5�%\��p1P�O�`~y��v��Wzb=�Cȕ��Ѷ)B��|~�����:*��޶Y��	!�o����ܐ���N7�����w�'��?���*)R���~�v�
�{��om�fR?�n����2�\���4o|֮��m�������]Xh	��̔ױfڢy�#�c�+�"��&AR��<�d!H���}:N8��o`@�@����}����5�q�QB'��b�/�����=�O��ݺcQ��I���^\p�M�+�Y�3��y\"�#5����4�Ja�/�pY�*�4���Te�m�_��d���X�z�=���kJ���-noВ�;p��6*{�i�ܲ��������>�����!sb���6��9 s����p���e�7�^��a�� ��d�� ��Q��:I�u�;���G��gP�$�x0�uP�����w����ް��g:�5����'�oN��T�P���P�1�	���lX�|k*����4�꜀�-���ˇ-% ������Y�l�;$'	<���-2��@���R���5�ګ��Lu���R`��[�w�Ҙ�Ys;��/4x�,�L���c�i���9TA����v�uo�e��&�]¸{���3xFa��^�l>���ۥJxiG��:�����u�1���)�W�ٳ�	،�����V�_�ڪ�l��PP�f�[$��{�<�~��m-@�*�ƈQ�K�O>����5�M9%�͒�t���ߖȸRQ�wJ1��Tj P��֭����r<�l��Sm�̮���=T���C�OYd0~I����Y�N� ��J���i<���s��҂p(R���<��m�+P�2�=�����1_@C��Ѣ\>��bd����ݿk���U�|_A���䎾O���g-�{Y窉B�(�h��ԭ�9��A��0s{�D(����b��&�lݢ�`���Eb��*��~�b(���W~�5�p"5����Q ���d:P�e� �����앨��sR$��L�^�f��Ӏ�5��.p��c��C�������������%``5�ѝ�'�M�g/��Yڰ{ׇ-Y��sdq�۾d�E���B/�I��o,�P+�m��40Y���[͵zX�FE#��g"c������{"Cy�q[c噥q�䢹s�7��ۈ�4�A(����	H <:���r�9��ְ�&M�Ѓ-.o	��i�Fc'���R!P�E���#���f��[������Ҝ�.1�}��僿	���I�~��S`s��p���?�^���\�FwFm¹�,^�BfT/��)
rV�I84�+��9�n�o)���)���q�#2��4M8S�m}_����ȝ��s������M�p���->|����M��ÓR���6�Iȕ���/���k@�qU���06Z8���}Rw���y��;�Y�EQ�af�\l ��K���m>AP�TΆ��2���d��}B��ڢ�8>������M2�_LsXD���ݦ�x;i��הݮ��b�b�u��$^����剜���Q"omI���J��s��(�q�菜��!��9��	��E�����k����ƍ.�A��x�J�,{ L��׽a��\{������#�Z�F󛉚s�6.��]�Ѽ��]+U����~�\�;
~�)������^t��<!���/��-mR�+P��?��gv��.�t�>�l;zA������8*��
~7Ƈ>�e1��Uk�c����K>�U+�M�ǣlT!4{p�&wU��r3af�=QHE��8�͆�:<gHS�q�t���(JGRh��	O\�Z!����>�H�>���R�1t����3>�؜�v+�"(�i��\=H�r�ڄ%��t|�y�����ܽ���zn���!l�x����kP\�U��8D���ʷG,�[���t��ۉ�����r�Jդ��j*�Ni.t��Y Œ�x��m�0�Ȇ�<�]k\�/�ӡ�+Z���Q���|���'��%�������_:��6��H�7����îx��t x�q�6��;�`r.Gi#�x�o�t��W�Tt��<X{!�D9x.{⇕(�ñ�Ibg�*�l�D�XN��Z��!w{����X
+�m�~ ��u�"s���y�\���@�`(�j�28�]�Ӭ׌y�?t���q�e�������M�?��X/��Z��l�|��ߌ�v/�]m���%/-��[�y��a�Fϴ�<SF��!ҍ�\�}Z|��Z��A��ad"�eT�Y�-j��!��olCn5����'v�QcDj��4�vI�,�#��Sv �k�8\k�	@a1X����-}�_�&)Ĵ�&?�յ��y���x=PWP�2�e�Lk��?�K/X�\�WɉlL�W��<,������S����Zl����^�hH�%�_rn}�����ڥ���`.D��!b��<�L�3�?X��dp�}D�bw`NU����:[}�_h��Y�����{��g4w�y;7��H[f�MN���2�%��M�Rx��%�d:�/���	�����&cxS��X�"�Y��/�Ii.�����mYO֯֟�C��qiz�B_*�L��4>~�g+�V��:��ݭ�|��_�y sY�E��y�0?�=j�l�(��wQ|q^�3(���ƓZ��k����;i���$1 4B&fK�LluX���M6�N���x�<ML�=F㑇�ݜշ�咶�)KJ'�e9�6�A��Rp��w.'�+���](l��.�Ff9�h�Ch4�퍝��,�����w]�R$�<���5ԕx]��N�r%�!�iE��d���B���6I�pf)�JJ�CQ��G�ѻ��^;��i$��KY��k�9�pm�7��VTYn��֢����l}�8��ȳ�Q)�s3S�x]k끅��`���Ӳ�#��UDMߛ:����J�� ��H��8���	P�f�{�8J9�c��&�~�ϱ�e�أ�f�l遜�U���z�1�����soo�MG�Q=�t� 3jXLw���>��ٮ8S���g�W!��媧��&y�Ȉ
oj�jN�����@q��xI�-�ʼ,~?׾Ǉ�g@�*��$@0�8������T{4�=�>���.�W���� n�x:E�`��K18�"��;��X�C�K���ݸ������?!�+_�(pw�o����G~Dc���<��ُc@t�����{x/�+�%�{��A\�T�M��R6�׬�~
��\�$k+Rhs��rylZZiθ�q���:����Jt�|rM� y�B�q܆V��Έ�q*4����B��ޯ-����"I�GN���m��bh�X�t㔻f�Xߑ�;L�s|)�!\��;
&��
j>�W5{L�/��1}c� !ls|̨xg������4SK2<���>��|�h��h�T&�����s{;f��?�=���`�e�[K_�9�U}����54�N���ܷ<�y��{OYn��Ԑ^��->H�?�<4G����Uvp)7�2S�%��MFR�U�­���U۝)5�xm��죚���e�h���/�W��2�o 9�S+r��i{CT���E	X�k'�������!+�p갴f���(��2�i�q��Њ/�x�*��kE��s-�+�Oܖ�A��l̺$���ˊw^'��CA�3����7qm��a�|�b���#j�ž�A`����І�bY�MQ��[����'*��[/s��45�ftPEO�����Att���p��f-��?���G�#/�Ly@F������e%���M�B�e�GpS��"����v�A��BRE�^AN�md�����X�%�I��sѬ�c�Ta�)���q*!8�;}}�W�TEv��gCs��B���\W*d���0D#pX'Ք����ىfN��`�}�}{��?�y�1�*��{�X�t��Wf��f5�4�K7D5��0����<�v�0@�?�-�!�e
(��q��:y������_]lUx糕K�@�:/�Yp��+����1��U�qT[������[����ֹO�Z�5�)3w�<��ɗ�B-d&�0���H��&�q�R� ���]� ��3�)!e���=~ZNQ��b��^�!��UfƎ���	V%�ݿpd�o�I`¶��W�½�P�z����G�rA��$B�����kU���sN�S��`�ʗzsS�L���~��5j��$\,�z /g��H������r�oEқ���*���|#9���%?۰л��sݍ��R��wu�����O4o�v�MH&3���[�M����"G���S&
� ����W:W����q�/{g�ߋ0�$T+��FqG4y�Վ�7�%�˧V��Rjiw���jh̩�.v��D� �W�q�MO,��f�ԥI���7x�2�<��	.}L���[ş^��X��z@ �Gk�P��((�#�A;.P׾8��*�fj���|�ni�*�$����cu)UA������<k������v�kܑr�D�����
���+m��J{���~�0���Sj%�5 �J����;@a��	Na�[�����b#�����\��0�]>��M�^#��m��|��|rC��6@I΁���{|��+a��	�<G��؁p�p"K���u�jEF�{��q�ޘe��"B�!�)cyvR4�|?5 �j���m�E�ic9}9�������Ј#��Sh��s��:G�\�_������"���;is	�g��T�����-hF}�*c��ܽ����YsVw�U��|�����{>���F�(Ĉ/,����=�X�A{�衉mu|�����v�9��.l��頒���lr��F�ئ�U\	�\�T�W������	I��%VR$���1�O6��j��'X���\/�8QRI�!WCʆ����V)8�vE��^_�y�#%O��L�-�)d�	~��L�-P�Y%I���x'���~q��[����d6�Gtf����& �;�,�3jY��$a���$��
XK��G_!g�A�2�c��P����W3��T��X�X��Z�J2�h���[�-j�J;@�����I��~��*����c��{���	�U������HK�f΂UU�B�a�yGr���a1�YĮ?"��~�Mb�>?�)`R�e�kdd�{$?�	q�]6��Z)�.%F��H"(����o��V�v�o���kW"�,u���R�Њ@ة�{f�*-[/���N�A�}��a���ۚ�-�Q�.�iE��QO2���'|�Fz��]��`\F>�o�( �����Ձ�<%!ε�t F��E�AE��.���#M!��PI��l�Ig�SX �W����D��`.-g!Vq��V��-��b�Z�R�ɐ��6��ԠG��g����5� �R����/�E�{�P�I���7ZM�6�XQSe�MH)�u�f���n�^����9��T���wBDeM�>�*�s>Bt"�ҡ�d=OtI��~����m�~�����0>�|2�K��nv'҆B�*�<�/���W��-�2L�@y�sF�0�}��I�+�f�v{�<�\P�(Z��4dO`ʺl,�)�V��W��rq�z1.-v��є�%����# �N����Ӹ�{񋙭��mJ�cq���'j�zR�
L��S�a��x��:�8�p����g֥f1��I�{4��}�u��.�{R���J�����B�NG���`�7���	Ɠ�(b
T��_�0V��㫨�ů����h���@�Mt�#��M�Q���@BTK�@�`a�"���;Wx`�ͪ���X�vm_�wd����+�s�=�����YALS�/D��˽�Vrkv�^�)��Kx���7�uY�4^{{{g^�sS�<�Os%+P���wbu��if4������T��}����r�e�S)|_HƠ&Vg���9(�&l�b��]�����UCc�Qg�?ҵ��/�k��P�'+K�J�*�;�����H�4�W�^�~#�ir�Fs�	j�=���DH̲2�,x�W�3���4��j���d(�;0�B���uΊ�_h���󸘿�b�M��)�a��a9�7�B�p֯	e/���"1B��ŕ�.5�g�]:���FQtYG
���4���JT%OºU�Y�T���d�L��V��P��͒����>;�qU����]�`+|u�H���gB����X��dvF9<�4��\�� JL[~��^�
r9�o�+�/�tӖ��[jj��k�l�e[~�|��.�삠��= ���w��&�%��F4�b�P���?�rI�2�/�T��f�[�N|gӞ�nZ�k���6��U�Cb�!�ԍ��j��W^�o�p��n��\���I9���9pZ���$ϊ 3�\:�:	����GKV+���Ny�ۥ_&����e=3F��/2����H
�/v��a��틔�ʌ�	dP�A���Qֽu�Q���EJ�����^�Q�K��髛6��xˆz��t������չP[>�q�p����d��?v֤�_��J����o����ͧ}�g�z�vd�$|�ō�B9;��6��h�O+��f�����fO����j͝�2úa7��$�����g�;�9~ɲ-�p-���ً
��H#�r�tY���
�c�9j�o��3�p�> �D��ܴVxr�K৹����ؙ8��DҌ��[�;��oJB��y^�P�/W��m���%�L��&񊫖)!��6�%��vԓJq|�0_JV�/A}z���$WLT?�VUH����>ɡ�R:4�ûX�Wg|����#$5u��>��`9��!	�_����$2��~��#a�U�r� ^��*1��B�'"��c�{!%viɟ�pЧT�	��k�9���.Һb�Ҁ��r�8��$�B��`_��U�0�e��l�!f&	�ֲ0��]A�$߯?@��i��!KR��j��E`�ll�ׇ@���s�\���������"U٘$�)S��TD[?W>��ߺ[�S�Z6�^��y����*���C6z�"82Fo�U��h��5�.ttqG6���`F�#F�A�j$��K���+)0܃
BZ >�L���jʖ�w�M>�=ܝR�(���m��R�d=�ޔ�4���������S2�4��5Zo��g�!�a��&���GW�G�g4�Z��7.��-�2,W��o��}����I"����Z ,�����A�������!Zԋ���1#�V�̏�,�;�W��t�<�bXIkhX�,Ԓ�� '�������шh�+��(�b@e��U/�f5ۇ�A47��Ԙ;��#����*Y�M��wl�i��3�R�w�j���R'L@<ŪV���`�b߈ǟAN�m��'Y�)�r�,*8L1��Q�]���M���,ȧ��:�&�d�&���oǑ��W?y�'�Ǟs���RF6���Fy����y3俊Ӛ}���X��4��v�g&����trtD;���V6oB�/2�|�\Bs �]DFX�ļx�I ���,�Fg�b*P1Ep���y_�t����a_��J���j���d��Yʑ�`̉G�Gz�/28�pSM-��2d�op�q�4���@2���5q�&�*�������Fԛ��d���rD�>\K�M%�r� �
}�,���vr��͉/������ba���= H�k�Uȱ�jy2<~�Q�IU7���b��С&&����V����:���
"��Cĭҙ��"���Zp���^���>�¶Kq�QzL;��{��tM��7���~�����_���Q��FH�}�+{7m�[��H�Ӷ���Z�$�Vd�r��c�:����b��E��$�z^�Ʌv�)��\|<Z4�/���O]���4�m���ԱFw�n�~���e��P���8�eTd/��Y��T 	��5�XKPM(~�jʎY�`��Yx�B�4��M��໸����:�묲�h�4��GJ��'a�ڏ�:�^\xL�"����"�PL�6hO��.��vг��#q^�Q٤q�%�����,��'�L9�s5|ޏ�ȕ���^9���W�XތS�gN������	���Zb����1Hꎣ�����Nt���*b�$%@e-�������M�:60m^$P�g�5Psa�sC ��n�Y��ۑo����\�Y)U�A2i�5����͌��=lv10{�ѻt��P���F�n���ȷ�`:���P���6���*j9�$�`@C�^P�̝i����x��S��:�!���c�-�h�>�4X��v�����,S�l�Tg���c�&qu�I��i\�[[�z��=Bl&L��_3��ueo���F��梀+)�&ʓ��Ϻ�L2�������-�b���8�&|�8)�~�E#_o�J?�z��nd��:/�ۭ�PH�2�0F�$�Z�8�N��F	�*"	��N��4:��չ?D?��1���!��9s��d�zlE��S���`�3�|�g]�,�c���ע�a檚����)�鈠^�����yi2�0�s�T;8�,�����^�vFe9���0��\^����aCYvыIˠ�j	�T�Q��w_ҩ=�W��A��ߪT�y�~���JkVr7����ZcZ~^:���9�(q�W]ay<��EV��'�s�^������SZ���oR��"p"؎P�@Z��,\$��+GŌ<�n
W�=%��W㿳��f����N��V��1�O�{��g�ĕ�K`,"ê4W�	�� �\~<�Zz���A�J�o�9첏M~&l�������^���};:���9�����8P�2����;��c5�yE'�������a�"��|'���7��Lx����*?2��BAXP��is�Kl+����N�ʮq�s��_]Q>R)�XL(�J	�~�¸'wl���'�Pt
�)�Zyջ&�����a��l@+���q4LI�04�����U�*!h.�@s%g��	�y!8':�1��?{�̂!����(��QV-6n��1�R�݅�:����Bƻ]�T�ܨJ������ݏ�J+f�ײsj"�vN-{�I�)rIF
+�&u���0�$����0l~��l�Jp/���9�������)ѫ(Y�u>,���G�l�qe!��2��A��t���v}㥴��Y.MSMY;o� ����Sh����}t�I̠̜��H�ȱ
G&�~�5;�S�K'�%U`0X����cs����u͖�qKmZ~�޵D�j�&�U]��T�(Z����FvxU��<C��+������U��6mV�B�X.g�"�^|Zk)0�r��٥�h���j���
$��W	��� ����"@F�����r[�}�r&���w}*���6֐���=��w�$��f;.n��KrPE���Џ"���>ޙk/�Y�Pc�ې����]B��p��:���{�q�%av���&�[���>GhL���?&��_���h��$�(.���yx,�ӓG�[j(�׵	䂉�S�� ٛC@2K�7o�
��'�舽�� �u���L��[2~cڧj�|�+
F�_�	�E��(���X�8ܴ_����� ��T��+���	#���O�m�x�%�7���&�ҏF7�)0A���o]��QB-W��A���?�6���䷹ W
�u&������.�]����]��|�>(0�5��W� Lo�d����'o��z�#��@񶚪I�gܨ�oÏ�d�\���F�����֮XW�*��3^�e�}�[A�-~8��y���9���Fl�NS��A��^NǪ[7`=Ȳ=u�,9��-/ܭ��Z�,�.��s�^�<�U[�������I�昬�򮥷����G4V�$�K9Ry�9��� �K2T��5]�6y���iZ#"�`���=�X��N�c.p�3�MV�r�|Ǥ t�鯼�toM����sE���o����O ��Dԝ!�M�ߏyD	̷��X�o�y� �g�q鿟�=<�>���r��5��"�s��f.�/�L$0m����o�[f�Ў�mfcg}͚�@�f��7��3�q�_�����YB�n�1i0��7�쳙�)$}�V4��,m�xf�-B?��oY�L|��}�)o�0�7�V`�ɞ���Q���Y��+�6./���j�._aXk�辰��>��ڿJź;i�A�����xk�s둢U�`?o#<Be�� ���f�­�U}���Ǣ.2�X��y��/����S0#c�����Ē	��ߍ��w4R���a6َ�����엌��]c�>j8�L�.@m������ka���J�ҵ��ٟ>�N8Ř����\�|�#MЀ~�O�j-��I(�!w��~��@$��J �qfCD	���t��o ��>�V�	����I���	��f:7�3�߉��
�1�^Ob��'=�ݕl��|P2|u;d{��x��xu{���x3�iFQO�#��_�	[��x%��+�����:��>܀�ɉ�m�]�x������XM�X'�E*V�s;�$��Q��W ��!+
�
n�^�D����7��!S�$d��Rj�P���A��vo�L��P�������#'��O�f�"�&ޏ3�L�\��B�N65Dv�k���c����H���%/\�[�(c _�g9�H�/�cd�
v���#(n��I[S��r[9�����~���z�vY�ʧ����k����-},���NG �i2݉�j|�\�#p�2�v�b��5*b4���.E�܌v�wJi>0�=�X!��Q,;"f�,)��H�S@U�`�@�`a��L-��:|"�" NG{�b�a�v�<K��[��7(�=ݻ6�G�$�M��͌�M�c"��˶���+T}d[�ڶb'4�� �cxee�S��e�YǦ�u�x���C�.�M5��t&E��$A{�;8��o��)%�~�"�$�$E��f#���*�!��k:G
^
�Ȩ�n��r;��;�����prY����.r�趙�U��s�X ���K��:.�v���U��#�bA�|f�{2��/�
���0+�ݚ >#��)�m�� ���2�%	���N�网c������[F�7T�9�C@�`�Ş�wT�u�	�T?q�F�y|�[0��6��8���ʋ�=�c<:}��O�9��}4���&����2���A�>��T ג/�y�`B6�M[�])��M�fB�(� ;�N?��8��)i�V�]l{�dk��|7Car�!σ��S#��t�j����* $~��{�����3�h&Ӂ&��Kɠ���<�^�g����`���/t��������Ζ^z���'���.��ɟ����L�*�ĉ����aË��c+爌V�)
�h���6�5�at��è���������1Y׹�un��� ÐeMr�,δ��+�h�E	��@鐫��|VD]��.X�͇lq��
x��#Wj�,	�^s��` �H49��6��@G�w?��q �x�9�{�����W9$��O][����Y������6ȇ�
�8�;�y}�B|�݉���D`"��� h�UU�Ɂ��+H6�7� ʰ���w<6��/V<���m5t/k��cq�T���H��a�XD]�S��Łp��O����N���n	ȿ�F�u�f���j�c����Zq��+rs�/��hW��ƪ}�X}9�*�n���ji3.>H�����h�1V��uG��(˥��l�Q۝�K����g��$/Դ�١ �Oq��o�=��T�$`��������3�Mu�6��J��A�#������R��̐�fr
vє����cQyӊ����Tu`�-�E�d����:p�apI�������>C�
��id�S��9ĺP}�I�(��jQ�Q���ma	���NY�I�x�g�B0�)��۪w��i�Я"c>�6�$g�����|��0u��,l�Ĉ �!%N#�U��nE܇z3W�ϡF�2�.HT}��{'v��E�ԫ��'+�� *(�G�M�iY��K������A<�,�&�oj�ã����5_�*����큳�=��@e�����ѹb���{ײ-�|c������P�@�]KW3�� 8)��UP}�W�t!{B��
���A�U*MZ���r�Ap��}�i�	�`Y�'=�N7�T^"nӚ=�MUW��X*	-p'Eg���G�]��hPkH�_�sc��g��(�"�k��^���Y	Pgt:���y̌ݍ�?�����b��/LJ4�,�ʠ,��!���af��0�u��}�Y�uÞ@WN�nX0��<ҡ� :�mX%���[�R�L���ռ.V��p�zP�X��D+�ڽ:�_l����
�G����x�$U�iMaP�p�s=bĻ��o��ѢlmO%<n�a�eD���a��2_cv�~ KȦA�d��+nzv�r��X�0��}��c�PuR�|~*�z��R��g^��<>�8Z�9
Խa3�S6$4y����p�ꃜ��	!�`c����D��,KxOf��緌a�������2��0�96{N��(��Κ(#�t�#u�uk�{�D�F���Q��n�n�	x�@r�Z�J��`,�oa$��E�)��Sm-En�>ś.��f��Bl�]�Aԅ(��������X0{$�r��\���+ۗ�+]1��m{R7�������Y��?p�:�_ΐ�D`yi��a.�����P3�sB���C�VQ�	@���P�Ȇd*� ��Q�v+�ZF�O�;���A�9�GA]�n�BwФ)k#�b���NA��y�:;��R��63�&���@�EM8�(�&t�7���R�ZbTv�(j��	F!<��>kT���qM��)e�ǻ�c�<��0�$���F1]^Z�#�O��#T�N ����+NG�������2�+���z�ߤ�,'l���W�Y}�b�F 1�����Vi\��m�lB����4��n�:Fv�|�|k6�Ѐ�| ��$�h���L��|�{�JZ��nh���ܹ�5#��ɷ��}K�᥾۵�i���K=g����h�'h�yWR�� �l�6�Spe��A�QI��~*�6�=��Z���8p������V)hwq7F��/��ܩܨP4�4��}BFV��f�Õ�
��IȐ[?e<l$�t7g�x�d=�N?����ϺS��"�hDnm�$N}1WH@D01~��/Z��G�a��@�hf���O~����^�=�Rz��zj����F�`�$*!3��)vF����L��ۣܭ>2xCl�*� �Ӆstl�T�0���=�^k�93�O!�dt�衈��J���{�;϶QgAm��+Qo0*:�8��g���Ȣ�2�ަ5G�OM&w��?L��y���>�eB�P]�pE���Љ��(�5����S��4�C���W|�3(�
<a1�T����~��)�1����غ<�[j,I3�*�G����=P>��9��0��CF�>О�͔��w�$��Z?�x�`H��Jo�E�T,�t�����u�ȋ.���#����������r���o6������w�g�����5�*]��BGn9feG����@�F������ޟ�Ǌg%����)����Ud
��Cg澌)+�DLS�,|1i�5`)E�?����#����g��zhϥ?���i}Qɖ�NᏦ���v��s��)O܄
q4����\�1�h��z-xwG;|4)�n��ynT�5��ᖺo�Y�zι<�,W*������*�eI���Fx��^�PR�Ipx�0�L��o�l�o�o^�:����<x���s�89Q/4vy
v�X<w�ebN�N�$R�e�Υj;����D��6%�c�kh8���G}u��P������k#���%��|Ydl�~��y��[p�[�(P�զ�Wu��{%~�^3!P���Qz�_c�5W:��Q�X�rn�c�����,0��u��	Gd�=�4�q$�rG���a2�zh]��Z1����1�f�U��^sN���`Ƈ�H$DS��9ю�d�����O�փ�N�ݺ�s�0�e��pV����Z
�;R�GͲ�i�@�68���9ɹm���7�?��&�%v,:ȫH�T�V��7#��K�~>Xm$)��0���L��+7���|P�X¾őIzCׄo���Ϡ��,�*>󉱸�����Ec3F/�;�4Q��M�N���������eN�ͨC����/H�eW�a|F����NT�����6����Q�ςؒr���f����><�J ��`��d8�?�^P�n0(����:�-\��,��l�x-�׏��[��1���ɇ����~���䵳0�-{�7�*�H�O��	��~�A�9�=����@ZZ�.H��������F��ͤz4*�����Ezb5�y0�H�j�ʚ(%�	�bnNU�5Y2��M�0?�5���J=m�+�NHL!����L17�{�s��=����^��z ��&7�*'�&�����f�cx��Y]��V��:ܓ�(vy��~���ͱ�>xD�@��P۩s	�>s��/f]�8�`G����ݘ�8m�L9k��孖�?t��ǼXg�������eE�{k#����o��[-��Ԧ5Q�a�ydO*��Z<xr?C���kJ�P�r �ç��M�|��fު���@�;���t[������9�ڹ5�[ŝ�%N(±"U�OT�G���(����D9���(Kc�sMgC�N#'�FB|�ZZJH97�V<�r=��g�n���س�BӮ(�9�Bh�_����v0Ѕ��X"/�K�5��)Òcj��ֳ�x�Y�[qK�ѡ��!9�-��]�^�UJʘ2(�vn��N�#Ň$�� ���-|V�s��:�o��
i�����3�L�[���C\u��B�_��������XEb�^��>_�`���9m�2H[���}�;j�	ꊐU��_�H�T�Z@t&ON���L��|�+��:muz+v��WS;�'��ӭD{g���:]S��1!��YK�N��Ə2�Q�<��`)��ެ{o���|؁e�c*w9��&h��FSr��s�=���C����j�ؽ��r	$���ۦ�'+��}+�Ui@����V�=]E�.��7��]�k��ǣr��J̯q<nW�ߩ�@q��3(9�h��]��Eed��N����u`sֹ�p1.jB����g�O<h-�����9�@\)�Ƕ9qe�Fܡ�e����C�������x����0��X�qg"��Mm��ɍo?�R
��&�܍�e)�)k�Aj�����c`\�S~�t"(����M��!<e3�"�8"���I����j�Y��˧�~��e�lUep����yc�ĩ/,��J��䕟n��ʹ-�i�b89�`��{�
&I�Jӝ��u��Ks�$�A8m����$E��_��Z0�qʱS�[(R��Š��:�l�7�\���Hy�0�[W����{J���A��	�ܰ0�YV�s�҂���ح߉vQ�ľ�y�̙ ���'��`o`�V>c��d4K�3kj��9$H�f������1BTı�Ӝ���<�Cٽ���Э�K�N��Q�C�z	е�OA��Ŧ�9�1��?HED{�'�N��n��s�R&/L�cr:��Q�Qq�?G��I>R��I��&C���CV;�7OY��.rG냹�R�G��� �j��������@�WVt�ϭo����Z����-f���'2�8��j�b�'�Vx0��h�<�O�m������R��X;aɑ#L�K�il�9�s���6m�"�S��I��V��)�X@���������|D��ej�t��i^�t�xb02�k�O�cuQ�~s���5k�&���9B�ŵ�+S�hoL}��	[�}.&8����&�hC,A>
�-醙Ľ��$�Ȃv�k��ŘB��������q󢆊_c_�Fq�RpGZ�i��*k˔�$ǽ�ѐ���7mM��҃���pS�W���}k��@��������+V��^�(�$�i1k0J3�ˁ�v��T^�����C��It��a�*��6Ц&�'�B_*t�2�t�i-�3��
ʤ�mNND�X�j�����V@l�	%��B&��p�a��`��H;��V��&SK�K�=���[֝p��rV{lF| �r�OC�8�
��0���ĉg�;��s'�
~��1%\�mē�M*�;=�N14�J�V��tr�$6R�7HgYC��#bĜ��)UH�(��~�G�[e�q����m�f��ŻH�/�{P?�%�'JF, �0ڧBI��h��[����-�(��m3ۑ�Q�G��}-��0i��#��&�}e{[ol��r��lu��֎L�|Y��k�Ŏ1��C��R���� 57Ǎt�������U3&ML�Jۼp��6����w���*�͖;�Nq�#
:�`�
�,�����>��x�������o��t1
�ǟ�"V�����М�>�<[��:����C-�}��&[��Vv��W�?�YF�G����H9(0e��0%��s~&�@/y*E�[��� S*E.�]Wf���=�l�Ro�(��T���M�\l�OM�;U�A㒈-�R�����ҴQg!i���^���~2�@��x�]�����������V�5���n�n`�7 j�e�N�@
@ �F#/2�$��%/��h1s�K1I�l�^�K���e�U�~f��ĸY!���S9:�[,1�5Z\���H�,�Ud\�+����J���0�^��>���9�S阷��ギ�	uP�U���X��&bX��7p��s�Z�L�N�>R5@	�-�핒7�{���A#w�Ǔ����0C�M0���&�_5tQi�r��ӽ��2��7�Y���y��wM1�a�h��.Q=��c�c�ʾ����쪃2�n'8�&ް"�TΌ�N��s�M�# �Շ�rA��3`�y򻲴���Y�E����랍X��PM��ضR�r�X��]&+5ڨ�d�jr��^�C�*�@���t[E\60170�KdH���pTU�M��T����3�q���R�M<�~��ۈ��8�[��,�#��Qm'��R�f�Q?)��ehV~xI��e`��ˌb���"�|�&��n�DhB��3�;��9�$����ј��=��F~���m_�v}��� :�QL��A)n�1� ���
�E�R����
Ưi��([S�`�j�Ҏ?�� P�0�:�׭=���e�'�v��m���;iO*����?�?h����!��OB��΢U�<Ή�m�9�-�sP˾
���17�o�����0r?�$�Fդ`<]+P��i��!K�3���`>���W�0;K	���"[�t�u�Eb�ut�F{������j-����0��l|Z�H��o@E׊)�͎6;�>P\!�M�p�&ǌ��F\8:��vʇ�}��۫Py%z6 �6!��/��#O0��5]j�"z��TeO��AWй�2�����k�lH�%"&dh9�6a�Q�����6���0������]�ć�n�#�uhF��{��㿿��qJif�`�l���� �Ѐ�Y�T��<��/��k�~+��W�ؠ*�h9�ξc�����Z�+���v���{���t����(�f�({TH��a�BK�_�`Pn��xw=
'w�0m��V>����\����!aE�s�"/ɬZ!�TE�N	�q���+@�xS�V��A4��fB�X&��-���G{��[Z4�Ɵ�ܱJܩ���P�Fk���fGٔ;�o|� ����@��_qݗ@�	<#����ǹ#"��"贛7]�˝�#���� !'j
��tkG핬V�mi ��`e�io������ T��/Ϳ�㐄�>)�G�8�]P�Mf~Eu%��X&>{CEL���\-�DU�]BuJc8�zvn1�A�Gd�̝����<�ir���AF�.�eeZ3����͢���JmSH+�'�ˌ��!���ycF�r�V��x9���J��;&�Y�0i�4�'����|�������q�[,`5�jPϻ���96��ߎx��o:~�~{��X� V��z��oﰙ:M�/IM����G�n�U�G��&�[.��A(V\��׳|'���o�:�-�y��p����դ�k�/]ڑ7�ZY��X�:�U8�����G��w 5��l�C���a���0>��H�Dk�&�T�ֺ����8��%s�h����&�q�����J̿=�:��&��rv~p����؄�q�P<!x��yF��t2�+�����r�vb\��2��e!��vz�_t����z�U?���������5�?��ќ�a�X�J� �+���%�;��O;���*���U ��E�d�oaဠ9�6�i"(��>�~�|v��ތy��/`��r��&@9 �d��7�y�Q�)���ҮM!k�ñ�b�ؖp9Z�������ǀ]���5�� J�Z�ZQ�����������P��I.�&y�IZ�{W�&����nNn��ehE��ӄ_G����^�b�����o�o�a���<Zȳ� ��C���"�އ�߱�/�3U�=f�-��uV��udm��^/_�6O7��qk�L���ߏV;_a;��A�c������]n�M;�Ğ;�J�m?�^l���#�h���Y��AB�S�P��,�2$�y���/�.��uT#e��E�'�eIY�o�.�����Q|N��M����Γ&Ȯ%�&�S�z=q�ym��%�s�ƙ2��������}~1���G(z�H�.���Et�7̽��#|!%������.�>����P�N���j�	�G`��[`��ޜ�Ŭ�ȼ�Y����Jě&�y@`?����/�5"�z���+��|l��}fj$~߹�nu����{�>xC��پdZ�A<c$���^ĤtCǸ@k�PB��0�:~y��s��ףVZG��-F��}�PL$פ��"}B��V�	"sz����dv����ѿL\�zEdֱş��x���Y[�t���WW�]+8�Q�H�MR%�n���p�AQ���eHt��O5йMKn�a�{��e0/j�����u�U�
������y�:��턕 �UUː$]J�)�2o ����%�e�gs�:,�	���ۺ��#��/d�J]z�P��*L�e���(?�Y;��V��n'��%Q�=��Z�?w<D�JSj(�?����G�ic��,c��%�;�_�׭�;KTh�}b������z��Uݿ�7?�93Q�����5�(]��y��.��0/ԴO������q�	�$�fp�|�*4�	J�T��eb��a�!>�EP.)'���ʀW���'��ز��
�=�.�.F!uJ�2�"s��*���Vt��dwZ���p�YpH���r6^�&ºU|�{HV��������ݠ��#"�ӝ��W���fO�5֯�Dh�z���_��&�{~�<�M�����JΠ鏟}�w��%��0��J"ӧx�>�J g�?f�aM��̓�1�2tv;�f�©�/� �`FQ�?��^qW(Ƥ�� -�����B�̷Ȟ�I~�b�:�KN��̢^��b1�Up����'�?ye���]�Z������߮>��h�״p�h!2�BĠ�'3V)�q��}�h�P;�k��ܦӥ�7����/��/���=���㉰��ɲ�H�Į���[C��������@��Q'A���벛�]���nIt�x/�iA0������F!�<��V,�.JO��Һ�G��!�
qc-��P�_�u_yO"-:�ZE�x-�L^�z9@�|�ƈ�1H�+11s���۞���[lN]�=��R����_f!u�}�+�Yɸ�5	�*([�Ե�`ՈmW��#��=�����>\�m��Իq^�֐�U��KZ���h��h�yU��k&BE�6��T���>?�%l8���N+V��v�̮Ԓ����3�<a5��fE�'6ZO�5ب�kE��w��#��N?+LxH 43�yb��)'Rt��v ���s�b���<M]���@�G�����G&�J�b3������0�ׄ�s_Rp��m�Z��xk��+��|!���/N�g_���*]+��}V�Z��6�׾Ή�e��1]�����\��������&�jd1A�Q��'�o�+�Y�E���W���CuZ��Ռ�����a�#�>�m�m��zwd8CE{sE�%̜?�Σ(T�5��=A�p�\Y�?\��%��z?����ȥ�no��z���1"	P"�fG�n��z�e��E�J��~�`�@t@o)�%MEw��[>ſ@veO��f<Qv1�P`|�N���=`� r/�����}3e�R�½ĥf.����|���J�L�(������z���Iғ[�H�,����S�'5Mx�\��ߙ��\���C�Ir|���.�����#��څ�����T���~�r�����ڒ4�dR#V���g�V�?�/h�7$|��cZ�tx�O,:4G���3C��23ѫ@yv	���Z�%��XJ��x.f_#�2jY���+'��͹���o,5G��a4�&�������E�kQ�5Z[��iw���-���e���]���<�P6]:�DU���]%�6qp���|�ۄ�� �T�E���ݦ:�`@-|�m�b�Rk���U�=��?$$�����gD�����i����U�X/�Ef�si�P��'���/C]�*Ψ�cv��|�p���ٲT���
E�$.����QX��=ej*�~�ѝ_��$�@QI��w��鼄H%�dw/bF�~o��x��'/�_��g��Zq�}���P1�"�����C�Z�c�ݔ����a¥Hʉ&[�W?�ȡ�1E-����|����w����{��J�oÀ?o�9X`�lU�r�R��*{�L��52rֳ�0��'��-퓬iBaW���;��)2�\l��nr5�_�h��ɲ����-j�2�%54��9��ϖ�ɰ���W�����5�^�N&��&G)�72�Sf��<������c��Bmy��+�g�d[c�X�F,�H+��	�y3��p�?�!�K��K��oM��Z_RKC�LF�7(��j$����V�⍓Sp���ϳ�ң��j��xE-�p>iʟhVNT�7�\��i�V����:��b��3S�g��P�XE H)tsRQC�$z�H��1Ԭ���|��(	LG!T������.��Z�@a���莻���T�~���竴f<E���±�>�j$r����H�?[U�/JY*�OH�����Pw@5�C�J�\5�1u��<%����2!e�7�~�&����	$��T;E�	�>�̰�i��u�����4�^h?i�	�fkc����PNE��vdI�v:�0�C�3"d��ȉ�f�߶���)�ǂU��60�M��%�"}eO�:E@��vM�g>����_�R�ׇʼr*>�M)'يnE3�,ˈ��w�R��:^�����J_,z}8���p��\�א�4D.D����,�{>:���:�c�[>����� h��x��G�Q�����u ��8�\�=�=����>��ĉ����ހY�bf.�&e0��2��\QGt�Ɠl��pa`����6�����*]2��a�9P�ֲE�N������:f�ahޝ���O6���)�a,��u$8��fk�.����cާAf�,8 JK�����Lh��+�{@X<��g�0y�_Qe�#=���������<����ӂ�?N�:��h�	B�w�z�ܢ�)�'�z�`~�H�S*�G��G��wI�T~��-��n~\��
�V` �\ο�:"B�Җ� sJhR`bU"ag�av�Ug��f ܮ8@�u)���!T�m㣛�y�����<��6����M��_k?��a8F]��J�*� C�A��$��S�N�Bk-כ��7/���wS���T��AN�uEp*�j�e�Mu=Ċ�~�c�޲�f�_E�7����t�Z�Nī���q?b�Da[�,�y�ߦَ#~���E幑�:6�g����gR .�5�����`?`�)0����Mg,��8~8��E��Zr�c��T';}��n�I�����0E�0M�/� /+mX� ���^U��������`��C(���Q��ב4�G��h0�!@��(5�&��~I�R鏾~��)�:��ي�As[<�
��t~(�S���ᗑ5+��l�_tRl��Z���S�`�Z#	���"S��o��]��F��^ �QF�YH�V4������>�w�6���˃,89ؑ=!h�����lo5�'��C(�d���oa���Yi�!�m�����U@R�f�4����y��bl�{�sC	��q�X@?z��=�|m���0"=S�s_��(l[�N���=�b*5^
�q)�]:�쇶��c2���Ia��Y�>�����4ͦw�U�1L��s��m\���G�n'9��0۾4�YLVT\�v�+>ԓ��f�U�[�[VMU��\(H;���h#YN��d_��R�)�^��C�K�|#<�_��g����6ծ�@�y�2�]^C3�)5+`[\������,�1���i���a{��d�����^Ϩ�����M=G��GQ"#^�\w��L�BN��0�p�f���G$�Mi���Q6Ĥ�?��=1����.EDe|���W�3{�R2a.���k[�W���Y��vW�.3ϐ���+PxJ�\^ o�Oŷ�3nͨ�K)O,�.��
͌�SK�"(�$�ݪ c3�n`�h�,,�#+6mͩ��Y;B+�	��$N��hh	A��-?pd�w��8=
��4s��B��HZ�1�P�!zr[�A����9��TPKF��T3Ҙ|~�{Ƭ2Q%r�m�y���)�ҋ�Ms�1Db�z�)�%��b��E�jg�ۃF�fs2�	��H(�{�Ռ�*�۫Z�͒�F+�`	O[!�,_P��Yc�Q�/qa�&�Ub���~�'��f+/�2K�-�;�SEO�x����mD�%Mz!3���C�:�6nx.c
�c"U~�B*�Q.�.�Kc"�!w?��I�N�{��=��2d�uA-wv���hH�@�-9���T���{���c%�f�W��gm��Vf�����)����qȃ�ߎ�����7�c�46�E;*#QَϞT2c��ĝ)�������f/@���q�Ta��R�f�_D��IRd�e8��9C�2�F�Ɋ;�u�b=�B��+�=�Mu9��D����PtXSu��Nvy�n�W��(�4���A�	�>��eh�5b�g�r�����eG�cbRai�9U!sEv�V��#@w���r�@�O�P��v���]�9�r�^{��O��X�� �C�˵b�(d�5��lQ�.,}8j5W}7���;7�:K)ߓ�nӞ�p��	۱&*t}���5�f8͞�-�L�y���!ۅm�&�^��V�������̇��o��wiKA/�����Fa��nLI�Ō�V�����:+b��E�q�._�V��}�ǵ3Zxi������[���ic���"�&/��|Tw^y� U-�I��˒�Yt��hf�ˬ\���;�H�4��f\�<`R���S����/V{C[0��˵F��;RÁMc�(/r��U�_��)��=�����_�Z��g��CeQ���� )�:��.��SJwS3�	� ���zB�оS��V��m�$~��1���-�@��.�w|��B��hr���'�6�x���І��ZS���@�c��ɿ��R����A�~G����I��-7N�F�:�ѪX"4�ĺEb��'��
������ue ':�w�=�#V� ȿSH�QYt��|�/5d�Tf�o��G�$�	ؽ5|�<���o���,]l:���==�w���Yno
�,j�|�ޮ��=�-�;���\��l����,�%�C^^)����d��#��u���^G�������QY�#{&P��]��pZ�%j��P�s���n
>����<�m��Ѿv���}�3})"����]�u%�|�Q�7��eVG�r5L��m�ȊK�w�c`�\}n�pw��7�����M	�WG/ �tQ{��4����H���u 8�D��9K��o�}�/��%��˚�^}��H�zzɤ������W���(]^�rm���}�,��@�`�H�3���Æ��?MBP�9��Cձu�鴤߳Ii�啝��(�l	Z@V�lR^)ǒ>�&F��RR�bjn5��R%,u����D�+�?���8\{:���G��`�9y/��G$�:M;i�7Jf��+z��p�������/F����ŵD���P����4m���G-o:�v�د8ߩq{WK�� ��/cn�Sp�S��y,z���$󃝳���kI���Q����Cg�]�z��HXYY��	�kQ<Qo|v�lj�ڿ�y�5��Rqy:
�dM���t�0Lj��z��ڷ�\�w&��tg��M��[�cQx�kV�K���e
�%�t�%>m-��˼Qn C--j���t�o��%���;�>9cŁ��I��@�XO~M" ~U���6&�њ�[���Ζ��^��4�T�e��M�0�E�����t�<��ׯ[�E�q�/K����⮽�����7����ӴR����>�&��jh�һdҌvm��sI�4d)�h�oǱvvn%>�S`J��I���e��%bS�Uʋ�t�5��R+�죞q���@�6/���d�����u�����ʙ`@鍇Q��
�|���Ü��)4UhI꾛Zv[^H&$O������+�a�ݬz����}���"�A�W�����+Zs�[䢉��o��g�����Q6��ܾ�>$W�s' E�2����ݺ�� *�� �L�:�
��ǃ6�"R��Y�c3�'���n�W�ú��j;�����z�������t�r�k�A���8ꈽ8�i-��-�r��Uj*]�����}Z�S�0��r��n����y���� l��W8*{�Q���u+�*����;��bgkqE��]���ܰ�ʆ+n"���=�y>����>��N�����*k@�H2�Ѐ�I�ڨ��;Ա��O﬎��Zȷ���l�+�'���8m�	��s�w����x^
�>��fj%c�5X�H֝�4�'����ٟk3�
d���w��^��\�(��j껅�z��L>������9�r�Ip�o?i&]�yi�������'�>̒�/7`�C�1�����Q\�(��~���4q6��X��ﴗZ^v%݀a�R"Ϲ�t`���'T߄��Y((L���Y:
�+���F�p�>\��a��}���G���>|>t
Hm�s�$jdP�w���,!��D/�P�L��,^<�=�%�{Wf�ǝ���t4�?�"hپ�U�H�s����]Z�Q˽n(��$��!����:
!!�����'�w�W�;�M��!�kZL{�=����� ��zz+3⫨����	��L�z�����۴.m�����<������9�z\$��1�D�8c��
�Y�"k�S-�{����h�,� b�{�C�v���i6f)ӎ%:nq�yU�8�X��Y�"_߮��#%��q��5/�\�0j�2�Q�/̼���]B�>�M��6�1.����#�DCAx�{y�t�Ko�9p�ˁj�e���' m%�|�8W:�QpD��gs�J��Ju�}R��l-o������W,":�	��`F��m�Xjk���hh�BbV��4��`D�ղLX�͑q�g��Iv���PdMݞ�6t�5wPbl���n=^��)��Nr`g�T?���y��?��Oa�!h6�°9P��͔�è�e��bj(�,@�����Hv�D�Nr\tj���\�L�9���І���y����&�A���[����8A�;zy�k[�Ѳ��A�D�(��N���"�SlA v��������>��j����u�]ha���
7��[�Ao❳6�~l���I��Kܗ7l��o �&�9B��XA ��9|������O��H�-a�Ep�,	a���h���1��E�ڝ����ޤ�F� l��b�o񮌉tq��6�w�PF�}��
��f�ߡ�KW ��� ��Ϭ�2[`�� �Ƃ�BH�0O��*bO5pIq��_mw8nl=���]����T��$�=�:�A���R"�wϝV�\C�������B.I^	ynU�DM ���ʽaX�af��$<u�}O���6`�:��`D���`!��\�z7�����E1=��	v�ވ+��7Y�cޯ)�B �00ڊ�t<��6&FX�.�]�Mj��>�IN҉`�M&��K��k�u���%q(��+�=�H>�#��H��G��ڣ�R��Mc�v���9n�����������Pm�aS]�#��]��Q�h�}<��[� �%��驯wЄ�l@�?m����l��v����"��דnn&<ٓFR�U'�ܡR�6"�"ߦ�ܦ�ǂzb:4�2_�s�%��z��R"Hkڷ�;��|��*��T<��{;r�\kZ#)8�����pY�Ջ�'\�bd�c�{�4�a�ݱU�Vc�8e#(�>��|AkJ|1z����C,q���FJ�h}�^G�g�0c~�ŕd]�h�����^NЈ;]�1����U���� �t�Έ�1xzl�M(�֊�AjIn�?�ݬU(��{=����]����(ټ��-Cf��M�VQ��W�/�TW;�Jۚ�{?�2�w�����oa=�v
p5z�_5
��B��s�P���hAw,;ͥ�Kd�
j���d�Z� �1����T�����F���0X� ���ХMdb݈�m�����S���Ā�C�y��E�镄�i��Q��i]��]�M�É��f�8�ܭ\��Qb�
7�'��T�e��7��<�7�Sˀ$dD�F{�f=�%uk��9w+Yo���S[���;W[]{F>x/�s��4���)*Q�STfגQ���$B<��.>3-�j!y.�W�Z����b�҈#����.v����!���tV�O񞥈ѩ���t$�����Ds���I"��p��@��7���1������ς)��*dI倣ӉD=G(܃K�7��;Vp�	��8F4Lq�6�٘K7d�a�~��f3⒰v��~��8�����o�+k��Jf����!���A�Ӹ��8��bΌ��kl�o�2�۝������m\�8	&�Ì����Dr!gHE�c�_L�hc?�=�����xᦝc�\
�!-�hh6�}ߛ�/�S �����>�m|�?��k^8�Y�uE�;��@�����(Jp����
�
g2���_����֡��ŹrP�vݣ����3���� ����G��2�"~U�D��ze�K) 9j��?��U��`(B�y�Ǧ��:
I�̶Uɛ ��e��c=,��ۃ�����+٥�YFf�a���

�~`r�f"�EmikN���Ɂ{��]�"�虸�� ���YK��Nr�(�}�Q���g>�
�b��-E��P����23cٙ+�UF�  �`~�Y��ӟ9�0�i�EA-%B;���8'���i3�)�ǟ��{!�������@T��oY2��� v��璮d�t*�~- S�����j��^��(>n;�jE�}`��,��(�zK�*s�9V�\j��)��ʚkQD4�#��1���|�Q���XS�;; o)Z��,�����X����Rц�#���5�ؖ��'e���J�ĩ���]4A�R������4�<á�sB�=���	&�lX��x � ��Y	�r����v���S�Rg%t�o�	B�5F�����m�Ζ�Ӎ�K�K��WJ\��q�R�T�Oz�5��vG�	/R�^ʗ1sg��xo	�M�;��љ��A�c�rz*�c��r�y�w���ƦP��@��o�кB%6ņ��q�������������Эg� �L�Z�=z�٭�����Ѳ�`��$0E�֏.�~�['[��>��yO�rB������aB��(� _l@�������RSڛC�v��5&l�ȅ<���c1�����mӜ��L�gx��t��0Y�q7��̪o�ƭ��}NC_��ƾZ�?��#���:�~�o
�X8��qm>Z�,��qD]3Q��r��x:L�|E�)to� n���r�ТG��ʫ���\F�XD���ߎ�̂�{��I�=�4��ul��C+�d�`�G��S�'T�}~+/l�W	ƴq履3�Վ���$�����'��޼'l�9Wo�/��w�F��ʐb�Ǫ�_���̨�x����UlAO�J���Q�����*��I���ǓV��;q)��ɘ�>�qt�{,n[�3+���׆��W�̹T�ܫD�ϣ���G�I���P� dKރ�r�mY�o}���,��r�s_5�;f���(L���m"N�}�;�(�L-�#$�Fp�'[6K�?� ������/��G��v���U�����+9Y�Wm[��]^�?^]ϨQX�sS��ŗ~p=�4�>W>��ڳ�b��:W�|��ޫ�9����>�(���~okDZ~}�P��w�!X�3pD��@����UW5_��/ZW܆�l�&𮄏��a%,�هr�r$ꛄ��B���C��[2�z��A�,Z��BĄ��� ېS$D�}��M��-}�_��Ҩ� 4�������J���0�}�X�w{�9�U����76�DD��E�8��J����1�J"��#/M6�U��F��T��Eӕ��-���t�&��;��yPT~����>��,}�-���m׺�eLѸ�k�7؄ �O�?����(;�!0Uu.;���K�{39@�V���sp����(ks�i��㼄��F"�ϱ1Ҥ�"e�<J�p��6��2O�h�ѐ�I�����Mk*�ae)���=m<�ȓ4T��$ ��݀��
���͹��������R]K�*)�eB�_iZ�1shNpf�aO�kek�ׂ�9j�y�%�#���"��$咾�^��\=>0K��,�^!�Y(Q��
������Fj�@5�Դ1�R���7��$nuE7]��lڌ�f\���za�O��,5	E)2�
��(���#�����Ϥ/��U	�3~Mo��w�*%3���#I� �_Mw$2�W�m��B�܅q�C��\������ ��X�k5�i��{ƛV�n c����� ��w��3S��4�m�,J����"D��;���U��tϚ&�)�Z$�Ȫ��kbM��г��^	$���-�j<+J)�s�/�p��k��^d5��{q��e�`���G�|�P��;�i�[���ﴸ v��^���^@p�۔��=>�$�]*\[3@r�����)4�w�",��A�3D��
��#0��f���1����M����D�v�'���B]b��.\')�����a����[�^0�nfʣ�M�����y��A�/�Bm��>�h��y�73�r�~�C��\��P���]�\
��PVW�C��/S����B`�;�����n"N��0iG"��7c>1 X��-�EFO� #9����<�
� �~�؉� VB���~ϕZ��i;������ ��Q�y����ϬTv3��ˏ��R�H�I'�bx=�h��WEb����{�@���y_@nc[�M�>���Ƀ� h���6���*�g�f���nA��鶛��y��A�4F��6�x��{9��z�7�f��:~M��D�Oc���L�S֙M����l%'��c6�Ʃ�]�;����s�7-v���L�qgx},�P��"�$�-�����Bҿ7ƞ�Wq��o|���y8�H���;X�)��A�$�N�AZ��a��>"��:7Bs1�=5�d�Zgv�������o9�URfk◽�n�O��t�[�v���XԜ=b^ίx�[�ْ���SL�[˜W�M������@���A����@xo�AI���x�z��y����4܅�0�r�h��~z�p�� {�Fv.�����k|B�o��nz�߱��Sȼd�Z��r�5�e$`���߱y/��C�$��gL��t���x���9�`�(uQτ��@��^�U7����F�Y<"�_<�В�C�?�;H���R
�~�2�W��kYp���d�ĝ�$��;8j��ӏ��X�M�����<L�����T���2�C�!��L@"�L�Sik�����U�uuിw����T��F��l�$����k!*����/%�w�Ȩ~���r�3D�u������a��1,�n���/�M#�yE���z�u8� � �ڌ�Q�	S�4��2�,��]L��T�	)�b��6*_皎a���ً���Ntx�۪�E�8��ye�\��۬;LL�i!�EB���kWEDZe�*�	4���͉R����/_v�]PM�{�w�T�N��G?����tQG��s����	Ÿ��~��mp��Irp1��'b]��r�g/��Uy�Ov�`O�*�RNuJk#�u6���Fǭ�Z4�Hcx���K�VZ8*�E��f]9�:H��}n�������_�.�_2�r!F�PL��\p:�X�s��.��RtX^�)w���T�+=L������15��|3_�:`I^5&:���7��`�ӳcה3�i#�Wp������_�w��N���v1�	��x����W]L��V8z`gH[�wZ��0z��zr���^��O�r���Vu��&ūd�"��������!�}��X�,��ʾ��F`���������d0
��{��߽��T������B$�4�뤄x嶔�@���c@4�g�?B� �^!�O�U���~�!�_6��:�|��&E��5MH�T�s�����O������E~'�'A5��{/4zo�KƓ������k�h�0��Tae��;N�}�0��6�T9j�E�ہ�ddePVB��.y��R�YbF���x��v :s�e�,ͦ�G�h��$"4>��گ��i���Y���@C�;(��i�ؖ�Y3c �?JBb�.�U�x�+WSZ�;�1�V��l�I���L�u;)�v�O�e��"]`ă��+@�p�]s� L6�8qv�4�	���t:����9�fK�;�3/��I$uڙ2x�i�=�����d:�N��#oc2N�SJ�M��Hᤘj��<t)1+*� ]�qu���Ey"aP��&��J����ڋg6�0
QxB�t�� r�I�����=�M(	mad����#�sE�W�2�9>�~���j��
��`��x�7�\��J/j������ū��*�GS�S82UR̍&d+�f�Տ�_��N��6*=q����h�5�%�T��(�Β.3e�K!�h7Vmu��31�O�B����*�HM�F��O�N�[+_�<htW97�by� F�^����&�=^�%b��g�w:?�u�7�[�#�S���Є�f�撨@��$z�y.�A6yV~�za�׍�S�k�g���3'�����ɢ�x!�#\�&]��Q��ؔƾ��w��{�+Fk�J���G�'���!"�UK����Ӧ>�I�^�H�e~P��:�*��2d˄�J���*1r}��������9���dW��B�4)���o�Ф���D�ͽ4?��(���5ߺ]���΅��\=x��Q�_ɮ�8����3̓��x�~��ӕ45Ɍ�Hw��pWO�x�0���Õ1���K9�m(�ە�층��D.��^Ɖb�n.O�?��|���</�,NF�.���OZ���kfj
��R9'��8����)(p�to���6gf�u�	�$�*��Й��rUڿ�B~�>f�=���(.�`$�a;؞�P�j�.�w%-��Kn��a��
@���Pe�3s�бzM�G{� �ߗ9揂B�>�BQ�(9���#��L��ʸ�J��0A�ۂI�g� ��Z��pXK4�J�&g1r�@ز��˃ +�s�ȼ�XF��x�]��1L`(�����&�� 6͗��j�c�<U��:�-��t��s>���o���W ۺ����jZ�[f�E�.��$逆����W��z�e$�pbW��9�%�#�]�˭v�^�ȃ�@��ݐ��Ad
[;�	R�dK�|�{�E�CnCcK����_0�n�oN��{�h�_�G���h{۝b��h^֌f��|0����ۏ:"#{�8�����1�	<bX�(12E<�m���5X�3Ú�#g(���vxky�On��˜���L���yWzg���ti"���q��(-d`�%-|�	ɠ�~���'���5���D�ʆ$�}�^e�%ݡ���ok~LI(����l�/6�Y������ʵ&R��=����y�1�������ϲ��V�Ż�����|��ꛮB�#GQ��	>ԉ��zO��]`~1D����Mh��(��Z��~��7��JB���'oO�.`ɭDԲ�f�?� ��
���n/��1��w��<2Mc`h�U��*�/�j��i,2�Z\�	l��ʤ�$r[��G��:�N)�4�%G���	K�Dr6��jE4V�/��i��>4VZ��"�: px��wݴ9�R�.��;�
a>o��x����g�i���7�Z����Y��sŁ�v��[���<.��^`>��?���L��)iW��bx�O쉮���^!����G�Z���fΞ�m����_}�S�.�R�X�0�0(�Y=�� R�<^R����0�����0��iֱ���N׸�c�	9cy>g�%J:��$��V��l;Jɢ�b�\�9��E�B��_𻮯0��3׎�[��T	��ٔ���
��i^� �����uu�m#��V��}�ICB��I���'��:=Q_�"&��w�f�#�iG� ��LŚZ����}� ~���@>C�u�Ri�lr ��� �n����0�'
�do�-�S��"M7�2[�ž�S�S� ��c��-.�aG�a�(��	��nd���D�b/S�k��~Ѧv/h_cy���齁tGZ��8s��������=f���[��{�f�9��C���r���	��M���9Tw���K�����(pzq_�y�|�c�8ܵ��\� �c�[�&���	�j;݋C��^R��_@�thr�M^�#OR������\�s���!�> p�z� �#=�>-�lwd�CO�&�+j6�10�ԣ< ��Ҋ����$�b떮�L
�[�H�<�l�i�P��gM��О#�E�ul��"�I埛#��ș�b�9>-� 	��%��|�{��U-q]*9L�x���A����m��h}-}�HjqA��T���wO������ý���8R_p��= b�԰|pXR�K{uې�5�4:n���\���1v�_c�/�,X���c�` �1f�_T_�ɤ�
�vDq�䛏��Гs���zUt���]F���.�2����M@������!���������s̍JH�E��x� FZ6� [;��^�;1�UyQ���M��n٪߾���mٗ9�4���xh���`%\�c̀�KS���Ɏ087�-Z�p(���'x�G�Ʈ��2  ������S�H�u��u( �u��G �˕e5YZm��Bgŷ��
�&��$S�����C�+���]�Im�7�`j)2�����d���� &Y��괳j��9��n{��&�E �tB�@�{���̶]C������Z�q_�i2��İǚ��AC�����(أ�h�����}�B�K�%&���4Bk;�R��%v�|Ά���U,}��u����K�v3؍J܏��n�II���b�iSk�lx��� =��H?� F>���*��>\�jzO�ë�9�"����LF���
�)������̫�T�a��Q���,�~u�s	���c�3� �")��V{���S7�ғ��٬!�o�"`��X��*[uv	�]�(�|��q2�}%wO�N�`܉�����3�\�%�-���e����1)��v��r�Y��Ds}R��$K���d)�̳�8;c��W_A�A%\%ʖg{�~l"wm�A��
��s����6H+�8�w *^?Ǌ"7Op� ��H�Q�d/b�<�$� ����`c�5VW��|�__1�i���L���yVm�}��	����A�c�ɪ�=��i=:�QQf�_P�ݚ�F���vW{Ұ1����h��}�TLC�S��#32�ǉ�8[}��j���ÚH�N*P�_i5_�����~k�K�����!�A��yB����%n���*l��CW-%�!��¤јf�r�/�d�WZ2H����U�߁��_���e�i���b?�ʊ�tv4%:]��S�,p�y'�݂-o��ac�T����-͞NIV!JF���Ԍ�uh��P/�
v,�)�6E"���'O�	K'���|����j��4@�}|.<����Ē:%X�C�4De��ٽ����)�	�َD�G#:���×F\m���O��l$\����/< f����nLϏ-8e��z6?
?� n�%�񠡚��������Ƴ�n3�f�7H��u����6�i�ʀ�
_�8��E�Y{,s3"7���ׂ��h���'B���4���{~{�٥��&`.��ĬV�����ݻ	`4���� �<l�y�J��~�?�1q�x����dj<��a��t�1���/�����Z���x�TA���j�T���2P Zh�zv�p~q�f�����J�ç��C<�Ud�̝t�œf�{O)�gf��իA/��j���� ؃
H��B�oCğ����Ǖ��^h�x.J��gN|��?�;�J�G7{�XK��&�n�;X�@)Tocζ��1_N��䰢2&�����F[w
���O�S�M�G^n ��N��`!�[��<A8B\�=nc��9!���9�S����[*�t#-�쌎��QJT�.6����^�#�ppX�7�A5v���"]�a"� D����0��&�y!�c�}��0�g��·*4@�f�B��R����W��(ʜ ��W�=6��c#�-�jzn�`j�۪�28��c��Mfþ��ɍ_3;A	_�OB�]=J��5�Eq�����:k4��n��d1�nnNu�v��(j�$A�����r�=�.��\�6��:�q�ް�����t��;��m5�a���E�%̣5����To�[`WԤ�b￾��"���3�Z7�ƌ�X5���f�b���j�
�Bn/T(�m��ح���צq���N�M�k*�O���Y��H�\��M��d~������������؈��='	�#r,�w室hS'�xz /�u�RH�\/w�R�
�c�_ZPYG9��OM�q�c� ��ï[��	�g?�л��3%r'5�;,�^�{�X��N#YM����:�VmfU����,�3��k{�zu^1Z���{������"Τ=��ͺ97�,J��\a���B*_�����It�� <Fw�G]�0l�����LG�����	���`��x�(	ޤ�={R��
�A��I���x>A_kv�.�������8+�����$��+�|
�ɻ[�*hN�ykzoJ� Krb�YU����K1\&�˳�Q�?���d���%��O�/m��e�+��������̆���5յ;N�T���^�L�߭;�HU>��gu��t�:��}i� ���]�0�E�������z��?ՠ���{�o<�U�H�y�x>c~�R����C���MP��/�B䆉{���	�_���hvLt�ݺ�(/���-��Ud�5���MG�Ͽ��m[T���3������.�U���P*4G�uRpވ���z�,Jc^uy�q���YHڪ.�(�#��ea��
/�Uq�k���?饌����N�kl�]tI�q�R�(i!"��ޙ��A�~�4��|w.Z����f}={����{"�#�;���k�@:=�j�������]㶵�2Y�/��Kl:vA`�r�,qҧ`�H��z}%uu���y ��5w�-;��l�I$0�À`��P�7}��y��Y�#��x�#���ъC�5�&�1	O�̿������_{�|`�"���E�zY}�D:E�{C W(w��ԗ� )+�F�{d[�e���K�}�6����F�x��}H����V4�&����N�kN��HC�Q���IШn�f7�)ABD��4�gH�S��Ͱ���D��o�T_$�*1>����ědѹ�����;6f��p�n��munF�c�+J�dq��f���Z<�� T��~v���]�����9�T?(:Qp�k�`�w� �'2�� CV]��n^E ~�PBB�#����5'X���sD����N��AHhc.���[o6� DvVݞz��z
���rH^|����_��j���8%F��?���q{i�y��>�r��D"�Ɂ��Pb��A\kRt�v%n�������׾LKW_y�#��F��
o!e��'�/�S72����)'�j�1IѮ%�+8cgb`Rp9��r��$=��}���cA�3瘟?��Cy���9MFB/�'ݖ6�����:*��H��;�M7�A�M`���:�`m$����ǔ�*���"xNXp	�d��)rq&r�%w�_� �I��|�h�c���:+�
 ElG.U5�͕BxM��!Ia�m$L�̈$J�]6�RÀD�+�=P�9�?�7����������2��ṕ7ů�Q� �G���tG?V��1ہ���d�����P��C�q��7p4�JU�[�-��'�vT1>���rpz^��nh�-v"����)����M����]])��&ڎ���K[���T�vu[���[�𺊦&���V�� pPY%7�ҹ�|�':�*e#��%~�R��x�]�佭aN��&�l��Kr��y �'	!�s;� ����(�� ��8���2����j�0M&>0���f���! �����c� z�Ȍ����Ϛ����|��;�{��G���6/��:��v�����q(� ��X!:�*D��Ee��� ���F��@k��S#�����(@4z�u�X i��ᾄ�L��4����O�yL�����OC����]�#����^�B?�`�O3�b��:��V_#�V��aR�=�GY��E45*I���-x����a^�Y����3:�dy�|��ƛ����ž���PF�^�^�b.��F�$���,��eN�ZQ?J����7ɨ`L�\O�\������~����aY��� ڬ�^�02r���y��c4�DagU���<&�.ػ�Z�*�v�M�SuB1��Mn8}g��8wF"˭��j�#$�MO�
d=���*�x݅�a4��myZg�u��d�J+*�ԛ[��:-��Bh	��ө���#�a�Fe�5��/1Z~��&B�������,?�)�/#��Q�\��&�*{�A�Zf����:X��/j��t`��K�B#g��&�Y�,���6�N�����,��P�,r��
��[ǒ>��ej}�Z��U��r����y|���\�9eL��6ǖΫ(e,�.k"c��3�E��q�`�Wa/�A���VܫWۮ_r+��Q�[(#�P�v�=J4��9f��C ���cb7��=�m=-08�
E|��'������Ҫ�l�vD��Ù�u�+�y�^mG,���_��9����J���em�h>* x(���MJ���pf�;Nl��k����ޚ�	�B+�T�� fq-�(і���y�:)/Ȍ��]`u~�W�D'��It���0>/4o��ɗ�>�u�F#/�'Rr��!p�^P1��g�=;�.��G�&�;![.�l��r;��=��y���,NrYx˰��ׂ6�_`�5�%��c���EėBqdj�V�F�s;Z�"��k���!"��l[�oK!�U��:+X	#��\�.���	�}:�m�P-B�7)P�_�Y�O>�e\nT���f<� `i��y-��ߘ6��FA4[-:Ɵ���窷�-(�<��23�4B7E>�\	��&� �/{�`}V�&y�tH�2��RS<8c��^/�`;:���*i�/N�I6O;ηZQ�T�"N�UQ���ϟ��m]�r��Q�ƥJn�:˄�ہ=��vQl�w�١?�.�f}�H)���6�#�dZi�Ih({!7���JJ�2���G���U���a ի������XZ<a�ո�����w�	�0(��y˵��B3���d�?3%� �}n�6�#����z�A��ކ��G2��o�^e^:GO��@�7�e)@�&NXK�����<
��p��#���85�6S��o
��'
4O��R�o���TdRc���4M]�Oo)��u�r�C�.�;&�a���k���Ovފ��X4,�&,�[=�ѽ=X���f7A>y���{U)�<����n4}ԗ򟢨+2`�I-,K�y�������2]ۯ��ʦ� ��a�V���s�.x�J���"R��!b�F�{N� 0��l�ta��z�W�E҇���!`a���9@�Z7H�Z��	���:.�~���>˲��/�[�aƵ3��QN�9j�c�{-N�;���:���'�A+�������o�pu	X8f����"��Л�P����be��v�p�Y���VE<��,-��+ �ʗ�R�2�c��-�pZ$w�v{hf�����Uɮ-5$%s�TNm��R���K1<Y�����d�P0m���4����j�8�UU�`<�g�X�ҙE#-�^16MNpdh3(� 3��f
O ���C�o[�h?���2s��tн#� �݅QB�Y�� >�}�y��U���t��=�"a+}"���m�;"�}J-�xls˳$�a�$�&����5��Z��+�F�[�-�[�j�7E�	��XeAf�4���d���-�~�3`���Ы�{������s�TCQ�?��� ~�R��S.<%�^V�и�@D;�"�,��-�*�bk�2�=�|8v���=�ھ�M�G臇2�6g� �8����r��yLFK�R
a�p�}f S4	�#|���7�����_��Vۯaq�o���5R�O�����B}��Q}�|�S"�:�� ��ߍ��Ho�:�7�x�S;�������*����B�ϢF����q�h�4����(�F��?�d�N�~�t�H�Cn��`5���]
��S��S��>u��5��=��OcD����!H�QfB<m���:Q�P��g������� g5�����0҅�rO��M�������J�͉�%��H@�?n�ɐL?�r�Z�˕�6�[�{ע��)e��C�$@����(��/|�<�r�֫E��"�.}��J|0,�����
ƺ��wq�^ǣo�����nO�G��ee�%�?��{��y�a���?8�4�Dq��-I;�d���������_B��5�7��
Oc���o;>����b�g�]R����
؊�ˊ�
6��J<1����]�F�Z�C4 �G罴���9�$H@��Z����o�V���H�Xds��Xq��������O�3d�(���<�iR��+����A`o׭	��  -`ѐ %����f,��ޅGR������i9�S��uD�X�|.8�려�[��kڔqW<��wm`a<�X/
��nd���!�U+��7+�X)��S�ua��R���*�xˡ�u�I5��9
=kc\����E"�h�)�<,-�l���,�P�R�����m�} ��*���=n��T����9�G8bG��"��:&�ظ;cr_=(�.�\(�t]Y��#�A\5�p�g�&NțY�b8#���1G��� �p�MUs���Ȁn���{�S�2�V�l'_L��^%�oy���_��[��ܜ���H��L2鄪Y~-�ˑ�Vr���[��mo��ֽ�2j��hT��c��J��&�s��8�%�g�$��dZ*sK�b�WY���Y���5��]��E�xzf�ۆ��r�8@=_f�]�	�<@%ei�j����� j��[�w(���QVX��@���w���S��s'k`�	��^Z��2�1���{3�ey�?��]��B�8�n̜/x�`(bi�Ly�G��ϩ0͎n�0���N�&s���Q����-wT�2���}|9��X�[*���BΑx2K�(��jj�ۻ{�� a�xdF��5��|�'�;%���-��_� 'xC;G2�n�a����=��o,2{�N1�(/s�n�u ����܃��S\�W��G�8V�Vܚ��6m�EC;�T�5��3�;0E$�n�F�*qP�w��>w|���t�:�,���
�徢��?�^�p]{���(Y'���Q�ijȴ��������|f�klB3�����מ1 ÄqDB������z�y(��_%�#��2k�{������e���ϞF0��l���%4X�I)!>��Sz�'���1�j;�-���+A����?L1��]K�zC��	�;}��D�cY�΂4�JI�C�� "5���pK�<b��4������R��ɶ��`H�Go|7�ν]����p��y��� �
Q͔zf7<f�i�
��6�K���WHW��j�>��ЂF���� ӌ[JT� �1���+�yb���NZ$Ç�mm[= ^�	r��7\�H4u�v�l�]�W����IH+b��ya��ƚ��]cX�Ֆ�U�Dct�LE;�P��Ϡ�o�Z�~붬���y��:(�i�qJ�k7�S)�X!��A4Tc�<)�����B8�R� 0$>l�[Ydax��5��aw��F}���gP�lw�-��ո�q|���z���Mx�6���^F@���,F���3#�D����B�+��wX+�qCn_1��H�gH2����0~��N�F�H������Q\������|�S�TΨN�H���:�յg;������P68�$N^Oɼ��f~��DψU�b�7^B/�l�e�8�?�ϳ歝fyZM�TĴ�2�	�������~k?<qH--CT}�9�Ybe��`XX^e!~6��_lጴSD5�d��R�~�O�Ԫj��a�ߟ�#y-��iz���9Dz�!c�.rq���%��ǟ��j�Y�+���%uқj3�yL8�Qb.��T�GLiߋ�9iPj:+˽ ��!~�W�m�{_����%��/B���Xz�K��̝�r#q�ѐXW�?�zEtSGvK�v�P	N�'�	�l��d��o��剰%�\�$����*�ey���������g'�	{����'+�ֳ4(�$��4BF�P_eqw��,�!�ڇ3�\��R�%r�;t� >,l�r�;�X��l���]j��Z��������v��Q��*a�5�=8�CM��^��
+�z���y��/)��e��^�k ^�-�}�}LXZ��w�h$�h5ؐi��2� ��$D��ʰ���s�5f�ѭsX<�t	_�"ʪC��5��B�`������5�2�|�%s>K3����	�e�bQ �F�m�!l�i~�s�.n��]�[�Ų�`TV�v7���݊/�;�	{��%�}�2ƣ��>�bp���0���[�d$���Bm&pfn�a��� �ݙ��<����s��q e�6�Z�����0������P�͑���c.�ǁ�*�L|�ŒXs�,�5mbW��o��0]ԘR�c��Bm ����6��f��+!���8J��#�d�ۋĬ�R���%}J�I�h�=�X�Xw��|W�0��0��e)T�x�"�n7r�EMH��7Y�~��
��K��B`a�'T��=���Y=��R4|u�&|@s���M���翎�91���f��Ց��&,gu�`�m�D�-�}�i���ǮW��$���
�vP�M��d)<m���3�Bkd���䌣1�>vB��G�l��ߛ,-<
�U��J�P-O?x1sDcp�ա�}�������m"?�1�Ι/��U"�ή(�ر)�s�P=6�a1���S�l�g�A���s�L��2+]�Ǆ�-͗c3��T><N�����듧����"�ӅA{L�4��1��R�жM���'Z���SʬV���\�%��tF$񚼲���\�����E��%Vw� ����y~3�;��p|�g�36 �۵Z�g�"���Uޑ�1�t��t�q�=t.�jwq;H����?�)X�F~ 0_�� p�M3L��u�����A\�҅V��2ԁbQ���Ye��1���1�s%�AݟX��~5M�kp�xq]w��^*��6���D�Qj^02,Ե����*�;7��m ���/�kI��)=~�!:�5��	�K)�3*�%�λ-w��c����W��q�P����҃�C�͖2EDO�d��钁�
���kM�\)�=��;�:9��|����7Gf�Z-�j�¾�$܄���{�	C��UO99�R���"�\] X
O�B
.��d �jj�έ��Lk���[*��c/h��������n��,�3����z`Q8���	a�7�.�5O���X[���r��婵g���!������t��8K��S��d��R?D+:u�	��%�K\�ʅ렕2W6#�ڥh�����H�����Ao�NM��=��k�t������q&1����a�|�0g��&Q�b�$�~�J�TvX�}4�K!�qz��	��qƻ�1jf�`S�a��6,T`�4�bb�C�^���
�X?,����)�z�L®o�v�.�H� �T8�yDi���C~wxk�P%�H���}N�& pJ��G��0�X�r~���c~�U��L�r�D��#�ig�����M8_r�	"����e:��=��Z������s��<���7��ܖ�!�|	�-+��-�f���b�Wݨ�<GMAԵ����G�zc�Ӗ{~�F�N��l��q-,��d�m��o1��D�����ʮ�LlH�;qBQ��`e�@�"@�>���ژ%��>��J��j�& \������Fj�Zz0kO6_ڸ� wJ��8$a�`-��w޾R�6	�����<�A��R� �3E;7����d�Y�8f���q��aL�y�f;�~���z����
H�"� čh�"(���%��w%�QT[!2��XqV;\VE_@���vvɒ�{^�Z�nWk!朸MʧZݥ:Y<�=9�'�O͸��ו8��7�|�jK�@��[�
'�_T�m��s�����z'*�8����]�oŁH�*f��:�>����;�:�)�Ȇ�s��͘U�5E�1�z�x�·0�i��U�w�]M\�Ew�ȕ��'gj0xH2L:�3^Q-ɱ
���NmaƛL���\�0{�H���*م�%�s���cާ�V���&d�l�:!R]���<�ow
��������,B�e��P9�WM���s�Z��Xʕ��#�@�Vΐ6V$����"*�N�f�@�B��Bs�� U	�8_aZ!���"aY<�K�s�aA:i��e�%�����ґ˭�J����7:Z��{�e�ܺA��W�$a���T���[Z1�o\��5��{okT��:�����A����1�,C��-������v������n� 	�JU?ø����>�!b?�4S+�A��b�|C���D	�����N�����6�|�.a�V�.�����Z�Z-���W�}����c���Zd��w�yNC[�����C�r�6>�,�P9�P���9#I� jEbJ�bH�<y� g�=�������j�/�LF��Y[|�k ���",Rd��H�C
J��q�^I��<W�����Es���z��zp�a~H��֏r��(\;��F�+��3-���T���k��,��'iR�%(�nd����٘*��}��ŏ$�xq��f-͎sv��+�TZ��ʽ�k�?��U\d� m��u͎MW,��b~�b	�⮖r,\~�32c�`2q�o�̞�R��z��񛗗�"`hU��=�"}Ӕ��s��R/��:^�ފ��}wC[��	=0�����}v��X���M>;�f�9�j�-�W:�'ͯ�+�!��/�[�ŀv���.\ʤ��P��>�G|3/$yu¥�J��M���OQ�x�������F������a�<��|a|	�6\���2ØJzS+�؟w���J=W�"�,
5��[~�M��Ǟ�����=�R)>N��.,L� ��|�}��N�Aϻw�o�����'2��h�eˡ�V�-��S����ѩ��+��v]����ʗ��NM|���Zn�u�=�+������@�C��3�T����W�D"-!
Bs��_�f��~!]]���6(ܦ����dzb��,K���P'JqX�����,��E�2i�|��g��Vmݡ�:�����3���
}^�~�����j��~e�C�	�'+L���;px�71Qm�<�	g訇O�7|��k�<z?}���oפ>��{n6E��+��]�5���v(9�6a�N��C#T��;f�*]��K��y9D�|��p�5��2(�\&�5�pcɤ������%gH"��(��њ!�����:�f �?.f#��jth���	+\:�"I02��L�}��F#\���>���u�,l�F{(�����X	�;�t};��i����~��*�vtS�w�Ϡ���O礝�D�������A�$�{QK���c�p���U֒1
�抈������,Y� F�r�s��P�$�u�U��V2�����mdRc�������t��ڱb�d
���߲�e��ovDi����JR�°/V>�..��$Y�)ت�����P��>7�㪧����۞K�5I,��v��ݩ��F��ka7��˨�-�� 8z�|�_�����0W���� �J�c}&�ipa�@�0����Scϰf���\�t���	���u�lkq
/f��>���9����I�j�U���ՐF	5BRoB�`��o6� 0�rzo�CZC�d�vS�9�����;�,)��F��lM$�0"�f��$w��y��d�W8�Aa�FF�ה�V�=ENm�Y��Y(���
Z��=�c�����ɧ�ߺ=s62�E���'��j���뎊���R�ǃ��u;Z�7�f���4	ުPʦ�G6x�ؔ�cD��ͼ{�kFv��y Ӧ'��.�Ө&��>��s��>{d���z���y?Sk�\�� ܱ.?s�4n��Rb:�yuH�]� ��ۻ���P %󁏯�F���"g�9̮
����P#7�nڰ/�`p�e�����>������Ѡv[�NG&N�k��ڲ�x��	m��_���c��%�;��w9�z%a����&�g&"�~���_����)��6b�IGW�Wb��l�@��Rk~t�4�}��bBA�Jm�P?E�X}F��j��ύ3����^U��4ht��J�:��+���ڵ%?R��']���i�����lGе��E�Fӌ]H8|��Ԑ�CO��E�L9�F��q��"������kB��>t	�H���_���LI�"�"8|�mE��ʙ�'��sa`Ez���(���'�!S�<�p�:!�b��QsF^�+%9�s�H
���PN�>�8l;�O�é�]�H�e�%�m
����L����s���wX����L6�r��3��c4��l�U�Ls�Y�uXk"�\Jyt����\����$��r�/�{�P�A�j�Wr[ލ�Pu�3h�$������}�E�E��(�B���Vc�@LЯ�E��3�}����Ţ>�*h��L�8�ley�俏�`�]�J0K���_}ὡ�`�gTe:Pq����{#��4wp���g�}bV�hHu���Y%}����j�69�E����v�g��Sb���eϚj���_X���-j���?����tL�Ys���4��(��$fcU�N��c��W�*��@�Ș-�/X7������u3b�.q7��S�OAK�bBq�̥��qN#���%-r�F�1J\9Rb�{{�_6�{L�ڝ'[��g���Rj���f̣L�ԵN����;d�f\c�=��|=J��v��	vD���xwK�T�S�c���A����=݋f�f�Y1e��҆f�^`4����`����E5��\����)�5��c��Vt��~�I9a��"��,���4;U������Cw
Is#�Ҵ@�ǈ�t�Ai�o�3�jiJ2G8:"9����/o�(������*v�%���P�6\��-z�	q��5���d��<'!���Kc<����E��>-j�&���<��t"F�0XeV����+�a��6- z���D?���d����Q��p�X��5�$�Q�,L�����Sۮ`]����g�|(?x�y<an�Л��мc�= "x��q��58�U�"��:Z~��6�����*�����X����2ǡd�%*�V�f�n���qr����K&-��>�k��<��c�	�ͥ�t��)	�o�����{��хq� ��v������������U%U��W]ƨbcXn�W��Uk���<�P`�7>�S�q�57bg�臂�����8k�����v֘�b M0$�!Pα���y|�r�n�z�T.�+H��ڦR�eɬ.V]���N�0�Mq��f z��\�������g����8�Y�#�ؗN��h�$�,��&y������<]ueG�vgj� ����7��>�����%7�+��5���^�(}7�����g��>�45n�L��ߍh�%�8(�@������C�I�����d.�����v�\i�+Vy���̶s��2�K��|uqG���PU��iM�I�Za$i_�re�kb'��&?f���:>��uz��PKt������Q|H�0� C�6�u��6y��ʶX���J/���ؗ�9Y%Z�E�~�WÅ��24�`��+�2jޮ���Q!7>hQrrFD�g�ꠑ��=�+�?���|�T�vn/���~���+)���P�c������1��q|��l��������ɚ���gy�$��f�I��l ���)aP��z+�:��w���a��~���h筷6����11�>��<}��66��q���N�J���+/9֝E�<K�Z�=�|ܥh"X��
�~�7�b��"��/C�te�1�����Z\�2b�\�cg���8u�;�g4���!�2�b�5��Аa���o�Ύب�$�)3�K>����ţՆ���o_�>H��[�ݮ� Y���d��Z�<�f���40���C���@R�Y ��8�>S4�Dj�Zߗytv$&��nDge���Y��PB)�n�=CT��ز�J�eX���u�IEc�a<6�!��K�se�,�мfF��ݘ�_��h�=H4/��S���t�r/���U�K�9s1��z�}_��Z��R$���b���.�g��:�#���V��4X��]Uk"�͗��u� QAX9|K*��zc���D����H^C��6b�����ɠB]rHD6�������O�,���3�V�����8�ߓ`�4�l{���*\>����R���� 9���'�Ÿ��g۴� ����?����N�Oۦ��x���@�A��=�a5�P��svG��V���2極q	����-1��qx���w�&��tػ��
����-��b�MY�h�G
e`�e�r`��h��f�\��~jJ<��c��q��B��'�(�V���
FWB�/���{Aw�u�{�ϴ��M�?�H:]��X�o%_~�j���������Ǧ��Kr�򪎲Ӯ�-|�vo׌��Z�O�@�ggۣ�P�:�T��f��kU�A�Ul��LO]��Ԟ�L�7��+ק�z�2�Z8�g���-��@ڣ�ֽ�HIo�$�����oqS5u�/yDlj�B2+r:�%��7g1S�*i/���6S��N�+�lxgY�Dŝ�zqG��s�|+4��\-�x}}��Q���o�%�� 1O~t�lt�65��ݪ�����|a�D�]ʷ���:)�`@�7y3g�#�Z����8(���;�:�^5��M��̕��bw�0�����'���]���S [�~~k�~�z�����k��I����D��z��!�P��d��1�U��=a�W���`�`�k���m)��<=]�p܅��Q��j�~)�x�1�mwߵ;�|�&�f�0_�T�[�ء�L�X�y���SU���f���ͣ��vmM8wh+��[�:��B�A�:�$=n\+��m`�U����_��k:5i���EB�����?%=0n��俸���Ke-��)��w��ˎ������~�c�r��H�7U�z�Qb�j��=��DG{�٪/�M�wj��#Ѯ�����g����-�L,�4��}LG��zqp`B`�\��m��0zF��N�:W>)*䫵��+��}���J+d<ȩB�q�y�_�R����8�5�O6��i�Q낍2�����5yw��k6)#�ъ���u�>��h�t|ڟ,���vJ��	^](
�d<����Zһ"�E�{������< �����[�xY+Qw��4��?�Ҟ��U�x��j2���w�����7�2�U��� ��U�âkl��P��;��&}8L��_]�2���#:T��Sy�Q18�6Ҕ��e!UVΉ>6�G6\����X�tm��^Z�&��ځ��.�x�8�.�Zq>.�i�v�*7c��Z�5�	�x�܄k�13�ɩD�{�<�r5��b��v��=�ue��X��tH�$u\P�"����q�����"4p��hp���	�O\P9���*�]�k����H�-:�8�pA
�3��@�r�KlYC �ay��9��Qw��6���
�(��ⱣV�=PB��4Իr��i�]��;K��M����v����΅~���[8�,�5�6m�|� �4�I�����,��2��Oㅐo|(�@7;�=W:oܙS�v��7��6���<ҵݪ�.��t-,p��$3��y80*��}8��3��>� ������ ���A���2�O�a!V�y��'U����r���WE�e��^�L��^��3R�%��Tr`�0���.z�(� ����r�Y��ƫ���D���G��3�d��nƃ�ÞA��S���z�<���O���E0m|j�N���hh-���,�P2�Z�=��M�.�XK�.��bǚΥ����X�u�y�˝=�\
��O��D����&�=Vr�}�(��~����H*r��x(4n��%{�ˤ����W��v����gU,��� LϧM�[�m�ލ'S� ?�,"�O2+��P�>��,�sV�����b�gc^��*�����m�J��>f25#sE��M�6ܾFz04��`�[�����Q1<��%�k���[3�ԯs}9���^8�0��[2꽎y����T�ke�d���R��,� ��M6@��lPf���"��Ɂ�\z�u�f�ݢ�\���+��&qb���<|�,���0k|��{�t��,kIJ��	�69&;�O�y���+7�V��$w͛rp�v�䋞�Bp�Ƹ���b�W����V����U]���Y~��=+qj,��V�O�F�n~��$@a {��>b&#���m.3��S|3�.�,�i=XK�(�4�	�,��x��*|;��i�v�8"��n�3�{��_���J��p�I��(x��E2;�D�O������d8Uְ�O�M��<�a�VM���s��3Ѡ+tOw��g���IԪ~@y"_�U��
VV���Q�ڨG"����e��;|��N��n!ȧ���¦
(�I�Cj��͹$µh��o��v�F
r��OR z������~���My(���b�SW��`������'f9�V�
�F\���F���IGz7�0��@�FN��(��Y^X�1��S1v�*����q���R6��i��f�fe	��-]`����H"ғj����t�HT�<�5�V� �we�Ju�m's�swB��|κ�86D���D�`Ut���G���M	z�m��y!��g��b6[放 Y��� �3�=��{����˳AL��/��PJ�ziG'�B��(0����F�6- ���'.i�ncOc:9��jZy�3̭Р��9�=ۣ�P�k+����_�|���@���7v<��'w������!Cu���Y�{	�������&6�Fg����r���.�*�'K�i�	�`�;XfBO�3.z�b0��@z��-ݙr�:a>����_��	/�>�rA��zd0� �,����P��~�wV�c��3\���(]&�u�\r�����pm���'%�Ǧ�wԐ���-,=�m�oi̔�6�|�砎���.���$I�Z���P�±�&ke˶˰:u���0�`X<����w�VJx���A�q�<�/�]&#�?z9׻V��j5�8*ʑ�Mu����Ob	M	c�?UJ~0���X�Q�����͚��;M�N �a"��u����d���F
TF�$l7 ׅ�m<'f����	��J����00�O���-h\{cB>��}�6�1�,���	���.j1�&Uy�?A�-�@�}��mw0�oJ"?�19^��DE^��g/&0G����Dpqv���l:X?�2u����걩�x�F����! ��1-	]��Q�ۃO��T&>G��	�h4�D�����f��.�ۣ��WJRp��V��Qɹ��v��nܗ^!��L5��#^�3 �T�i�J�K�q3�z�8������;�:!�l�I5��y*���Dí�����k�x�����Db$	�h�ѣ�������#�2�?�p[�B�ʶ��)ȸ++I���:3Dѱ��y�:H����U�x�5��,K�̵6��7��O�cSo/���!s'�����w����c3E./k���d���B���e?x�a _a��V���������#?��]�lL	1|�Z��B#����)�+��n�5Co�]]��t��ޝ"�uuE�k���@j���AϦ�%
b�S�M9х!�4	�E ��T�D�@�$�I�:b���;.ʜ�6�d%@!��c�]�W���;L��P�u;�����в$�P�~�&����[v�%N���f��i�ܲ�^�9.p��X|ܔ�/*֜�����ڪզ�T�>-l7)պa�x���X��`�2�%"�b�<cZٗ��,�����6ᩥRϴ^����/�H����W@=E��?N������p�}�N�=�K����U��6B��ړ)�T�tԲC�f�C�Ot���U%s�G��)Gb�! H|��4{֢[��w����ʓ2�g	��=��>,g.�$�'��q^k|�>�O�g�H����e*׌���;�"�������dThN��?(i����6�ND�����M�P;n�}j>on�\�]�>g���»D��{����L`S�]ǩ���E<^4���H���c��%v�g��EZ�ICf ?0��	`v@	��,��5}��!�p����)9���T��5��M}�G(�T�uFP𬛮���t�ŭe��
 X�U1��+��0 ��Oj�[g4_��@�a���j|�I��x�Qf=Ū���-����D.���e��~-��Hă0@6֫^ۺ[��d���q)���q���X��aöс������P�3�ډ?���)�*H��y��Le��?=V�p�ꞜI.���� ��.�'ݳy��a���BB�$ܻ�'�&hA��O+�����Y'��4�y�u�ZU�_1�;4������ވz�2u� ����~�goH�$��a��B���6o���\x�r=�RM|�!���(�i����C�\9:�;���|���?o���:]���Y�X�5���P(���� �&e���6㨥䪥͕��|�-C�v�k��+�#�Q;5�l]���ڮi+G��kɰ�ؖj����#(<�C����H*�/G/�OZ?R�#���\s>�E\�U�_tp<���9 �U�ǵL��c�xV��0��ւ��bHC�uny!����B=c��zʵ=�Kj@1�˫���]O��3�qr� ��베���&�6!X�H���W��[�!&�h�ǔ=L�B��l�'�*��M[<7��A,Mh>tq��>�̸"��p�����BsDSᬥ1�3P�:�[�4���f�7b��GIW�a�b�Qh[Y2�Ǘ� @�R.x�^��~*m�+�C���O�|{mᾒ�|A�yni�a�F�9���T6юb�ܞ2�:�
�8�s�1�>b��y8QhYkk�h��ql���ە���q�C�|h�"�c��s�@ſr�u�%M �w���������`H�I���С���dZ{�n�B���g�&����4�6��<�����	�-�*0|g@V�ԵŢ�ցm�}T�c~��Y{����GsC4�=C������*S�eqX��~�vK5�׼n���Ո��e�"��l��W����/8�C(��������
�x/��4kSP)�i�/�t�|�1��.��%ݼ��F��Z�??>���k)���k�����D�N(v��J����E�a2�2y(�Q]�g�R�;�?���6�b+�������h��� �Q��X���pU�X+i8
 ��*�Ҿ�X	�V��D9���U�DJ�T�B�(��ge�����ම��GG5��h�I�j�>���Z�t��}L5��t/�{^(F�!=�M `�����6�e]+
���q�MA�Li��t�=��59b#�o�rPO�NPc�h\�A�kK)�MU^����R㻺�����9�eB�쐓�k%2V+��B�$��E�X{�Dpg����*���x�@�X��Y�_��k����y��R���p�A.T\��p����A}�91!c����x�{��b��u���}=)��Z�4��ҭH�̕uJ��U#�|�^��l4�"�8�<6J�xzł;x:]Ji ��eǓ��[K�:���l{>��G��a �#��@~�&�0fhhg��� ���6�TJ�w��U:k�o~���]�����"v行L 3܏�r��п��{�a�keرך�������� T=y��2e]"�I��0&���?%�X�2/�-_����_�g�&O���۠�gdt�9�iVJReT�����s��6ghY��d]+���3<~F�����Q��\ڜr�N��P\ �rV}��#�`�'_v(3�p,��{���T|m��O
���D�X�+�7�%;pQ*g8�$��)�CŜ����� �2E�m<��,����h:����l�J�9I���Js�O�M 2�'�U�1+����3��L��ˢO�\�b0�M��=��gP&]���pݳ�	�?��{�TE��m� �,�Oِ����p!��'�9��?��ed��g@�����N�G����Z�~�9�qܠl��e	)L���Y=2yԢ(w���I�[�0��?"Bj���u�i��o{�W���a����L���D:ة�����*ǭ�o{7�zr�/8��މ�x�C�<���H|L��A�����m�u�Z�r�á�p��.��廤~�X��VC���oř*FT�t3�jf����*a�N��1�:��k��9�N?�\d ����R��!ߴ�U�Z�7�����fXg�q#Dv����H����8.>��ZC��[B�8�j֛���1b_�s��k0?�k����n�=���hJX�uS�f��L���z�����ՂO�W��11��� I�/����k�_bfK[�[�K������� �:���v��Q�����s�0�6~��@.T��Ŭ���Kc���Ҵ���9ŉD��0���:/^I�78�U��R;�_����r^<��򟅉��R\ڊ{@S�<��P�"o(敫B������aA��e&��L� =
�Q���ڄ��Lꈗ�󠷊~�-'eW�P���|� �[���c6�^�ڊi�ە�+ˍ��PP�<���Ō�_��QO�('����i��d��es�=C�|������N������#s�<`�%��E���;�J�\HXH}y��ѳl��	���S	���]�x.Uܽ��� ,���A�8���0�Au�<)��O�ʃ�:i�`1�k0��a�\�~���"j6S�����*E3?L�qT�F�&�,��ƺ,n���%�����R�8�i�prH��u�^�� ڇ��i�n�`���Q��5H����0�P��������讖7���wl�/�pV2H�]�r	��Wk���i"�:����[a�ܲvj�y-a��4�P��\�62=��a����t	֔	�9��^�Y��\�+yb���dR3y�z�]��T'�Hi�n�����D=p��+�U0�-\'�x�#Q��fsY~�u`�7i�T�Px���7��5<
����Z������t���NR���y�ǙW�Ay��#sp��Y�_O����@��P����r&-f�;�F��
g[i��H|��?��z��U����9B���D��3A�nˋ�@��>g�7�p��
ڶCB�����(�?�_���TF�Da�,�tJꌐB�e�.u�� Z�ďfՑ��%�N��lL�8F��g!���ﬕM�Tm��#���@b�N�SF\���J�q��S����9������H��U���ďv�M��}���`S��]G[)T���z��-��A����nF��\�`�$E�MSMu/�D�V��U��^X���'��ݨzk��j��2�gٙ$3$�a��J-:<�^[���j��m��z=��䨬9�w�kA�:��\������nd���c�6P�$��P�+ay�ve�>�����l�q޸O�w�C�8����e��ғ.I�4!����x�r�!�#�#T���*L+P��~�5��85�e�c���W1�}���<9(z.i�lC.�#�kZ/JvRb��6b�
����4���x�F����a�ɡ}9��1���'7�!�j����e���]́lf��=���A�[+m� ���s�fR�Ҝ9�k����l�y��A�f-1����ݕ|��$�_S�/���k���g������D��u�l���}T�b��	�Cv�a=� ��p�>b�ʈ&N+"nSoݍb��^��HP�w���aM�U��I������:6���,��w���P,M���N�,��o�'l����AM���9Q�fq�Z�ͽ�ڭ� {��]��(�[���Kx��G�13Jv�����q��K�;�9���E]ɮn625(z����\J��,d}�.N�a�q<��0��[�;!8u�7��/���J:�\Spҿ�{�(N���Th��VV��Y�7���� ms���uBҚ���<�O!�h4�)��'�%�B������s��4v�t�t�M�� ���$�D��i��iul\+��=<���F�U�C #��A�S^`L��n�ٙ�&��9��nKߦ:}�>�����o�̐�&��*�L܃Y~J8��]f���D���������$+��wtw�߿T�Y@Wsk6�H�4�m|��2l竢y��Z�X��g����ީܭ+�(�0]��͐m�!mrz�+3,�s�^;��;{�X�D3`��Z�S�����B!��N=Y{�u�nzF9j
K�8�Z����t��h�x�VfYGD�+�̨��%�o�����(�C���1���+ڥ����<}�ɂ̊�ڼ�f��'u	�+��̿v�i�?&��=��(�0��c����V74��C��l����y�Pbm�sd�¶=�u�n	��-	*�t\o�p�{��}&Z�0�� ���)e��yq��a�Q�6]׎�����F��0���C�O��)R�j�ڎ�������º2;���\�P�1k&�cn7�.H4���I]�ng�; q�Du�ӭh,�K��M.C���½��́C�wFw��r"���[=F6R��m��[B�܆C��������������L�g(.�S¿#p:�E�M"/JG�I28���+oU4�wr���}���J���K絈&~[:B�!ִ<R�	���XqNr1����lG�Uu���܍�!Y�
>��_����'y ��f��p|�
�d�d��=3ZS.�刿֊��˔a}L�B�5b$��}���͌}H��5O ZPػ��G�����r�]������ �ȍ}�w-b��@�an�:�x�X��e�:���Oj�'�V�_��ki���Y+Ę���R����%~%�����r�-���p�/|�i�L�oZ�}ug�o��Ǖ�z��d��(��%��� ���Y�G�h�[����zG5w���1(h�\P �p)A��C� ��~�5O����M�������@�|t'���z���T���Ts���R�n��.�U+Y�%'�@I4���C?�#w%�B6b�Y��ә5.cƈ�_�������͠G��U���b�n�M(f��������g}$4����hUh�o��vQgx���q '�w�QPq$5$Y1;���a�l3��� qt:���4襅��a$I��"�s�1@W>�5�n`��`�iD(�3���p6J+�`!l�A�Z
8uUK�x�������[���n@�Q�{��*#'4fH��t��}�|�8���r�C.(�J�����]?3�֡���j�[1�=�b Wc}s����!�z#"&����u 3@�֎Cz���fzlll��EW�y�Ǟ��م��K�R�
n��)��Y��i9�w\�ᙠϪ��@"`�80�w�v�I��vm]��%���S>�{y�1!���Eh2�1����l^ۃWe�p{!�Ű��V��7$ʕ��X����@@3%������Ϣ��Kux[+ʼ|DC=��Ӭ�8Apqt����$�I
MV�g�찮�'cĶ�rm;~��s���fK���$��g��D�fV|=g�L��V����D��\������3��5jɲ��j�}��PF�t���]l�~�Z �+�Of��Sm��&n*ɷg|އϻi��rgF~��I�r�?6�{�Մ�(`��yXɋ?�ko�G�(/}_A9�,r:��+�>T����˙�%m˛�͡�گ �]�\���Z]<����WY9�O���%iqa��{��8������۟9�u��3��9��r%λ����\|������������C�C����'x�x�<���:��cG�y���#��ʨ*(CEI���T���y��	��?�, 6NpF*�j�Q[��q������UGט�a �fXj��j[�Tَ�c�����j*��i�o�����W;��3�  GI��R;��Uñ�9y^~��*�*B�j���'&�gp�����L;�Dʭ-D*F�S�n$�5�*H�f���1�n��gmj��i��d*�8�2�t�A�3���g��Rt%�7���ÜGȥ�@&���zs>�8���0���������i�#�����og�rR��tݜ��w`��d}��ռ�=�<���7��FE��[�je��ߤ��q������bx0�ۉ�pۑ�4�CR�����C���VTo���:�ϧ�Q b�2�S�-%+m���2���ރP�ERs� L��Ju�%��dD�6�ZFH��P(�fR�"�M��"�$
%%���c��"��#/`������8����Qy	Գ� �[qc��&�Y�,&r�5G �_��nN-��s��V�B���'�>)�u��z^�Fc~�n��j~�/s�2%�y?s�=(E�P�|뒞P��yr�:L�|�K�� >A���D:���e���p�#s'�ߟ��F�c)?��#��ǯT*��cwv���2m�ס�� �M�o3C_����%Gⲝ�1����В�w�¬���ܙ����^�>Է ���	����('5��#oh���L?n��s+rǰP.7�߱�<��J�z_'����r*6�zi�L�VeXbA��Lo�)�#uɾW7Kl��������B��S���L����S�'ϑ���X�Fx�a����!.�7�3�*�_�-Vo�tK$M�V@��.���s'%$U�ʂ�'ȥ8�ۭ�ƃBD���#I�_I�LwdA!ݷ��� ؅0�]��E�~c�E@wcԝ�����ة�n�'��ɤx�b�͟]����k���2����%Ѿ�+\�.�R�O�7����c���X:#��A�zT����S��1!r>9��K@fl��Cm@�_������x�CwE4����H��]
��.�d�� �E0*�0�x��/O����:|���	��D�]c��0��u�s���L'�}������2U$)p:�f� �(��$~uʏ��dH�9 2x�c��[δ��Qr�g؜G��uH��r�P���J�/:py��4r������`�ԋ�/ɀ����!*��RZG]O� �� z��۩��s�8S�!gB��J'��� �e集k���$)�k���S��K��U=�v`[\1�	aɂ���>r�)p�V@��ڸ��r�̀ZQ�������W%����
m��Vt�dH
~G�۸8쳙��KvC×
Iz� ���D��W#�r���s���O����mW�QE<�A�z7V�vǴP<Y@d���ϒW���f�N\ Z�k��^��_2	�>� �E-�����u���AXǙ�BX�%Y��a�G��0&l���3��2$��2B�Z�ZԨ0��C��|��cVL���˒��M �T�k���@V@K	��' ��{�G?���ډ"Cz"M����Gȓ"k��0�'J=q0a�.b��k�&�G`z����ӱ�N�\�򠅯������M݇�:}*�����e	�R��D�$�+�qk�RFj��Q���{.vxƛ �S{&�_�zC���N�p�E�zd�Z����C<A�}�a"8�B<��k�:�]7�v�!�h��w�޳$0H[uuƃQ�hP��I����C\<[�<ݮ�C�{%J�x��1D!ID�� '�mʌVM��v��Ԋ��X�i��w$;3v�KH��C@�oâR���(^�+��""����oc��%�4V��6Ƶٛ��F�r"��4dt�����EKb�f�����v9	��oҙ�hI����c�Z�f�z�G��\0?�U��mQ�W-��֓T��&U=�l��j��$fD�}�yt�+��mllvw���u��NSp��7��ƽc<_���,��L��L,!@�����z�Fp��Xujd ��pG�v(�C�e�k[���[N} ���Yy�)<�*�	�����gȽz�	i�uc���2̩���K.�����
�f��T�����kg�P���G��c����^���/+�Mr���T�T��ͦ�|�ܰ,:vԧJ#�	;\��\E�z)����rU��V�׼�VVFÀ	?e��8���ǝn
�s��tҪ�2͙�O���N�X���e�HSg�f^�$:�љ�]���,"=(��`�o�O�P����`� f��.4����M�*,��c	��'�X�c���b�ѐ��8���a��+�V�q�ؓn�2�Qj�j9)r?}�����~�SXͻ��nG���b�m-/	��8FM�_*�t�rw��zmZ*`��X MG_յMO`oi��a;v�Y)���pj�����X�5E�]��E,��G��ܵ:E�$�4��g�6���9:��2�S]J�"�ߤr�M#cw�QY�$vtZ�@��T�9��Ѷ���nq�1���HA���"c�,�Fٿ����i3YŸ��3}�Ά��~���uOK�=� bc�tk�~L�i�׃X*R����C?��ۊ7�P�ځ%-j���يon�P,迁�纮u+-`�?�%/g�ޗ|��E�#�pj����?�b^��{�����*�i!B,��Ӭe�	A�x�S�K�� <����S4G�y��|��m5�Z�|c��}�n.(\�����l��}Z��1�>�o2�
�Ɛ
�,�Զ�TIl�m�{kqL�G��?1���~�lw�˿��;Ҩ�N<��{̦]��t�_��m�{'d3E�Y�V6���,�Z*�ð�V&'��4sQ��N��B�wi�,�X���I+R)������$��Vɚ�)���6λ�K ��3��q߻.+�^_��*S���V�ub�상=r ���N�	��Ԛg�|5��-|��-R�ΙL�Ax̑���m��e��m���q��s�b��l�k]�~�����@Mz���� Z�K��f���1E`����c��)pp�'��'�U�m���(���R?ُ�U�ž8`e��Pk\����Q-�OI�ۊ��O������'c&��3��� ����\�����x�&��<�ϹՍ�>�
"��=�g�υ1���p?�_��o!QU�W��^Ϯ$_r\w���X㵔���nn�
ʧn�h
�*��v�ҜFĿw(�!2A0c�ӂ�!�A&�w��-����pXg|K0%p[oʘ�(�I^�$�.ƣ���8�V����(�(�!\��tWނ:���h�O�
�pV������MΎ��x��$� g���e 9��j�°�SH�KKD��X��.$�|����$�N��� u	�,I�($����1-�Z��������8��ͣd�eeh�:�����B ùJ@��ۢ�Ӈ�G��=٭��K\�,%cl] 
 �$�]��	+�&A#I��c�I͜w,ـ���� i"����� �G��73M�j��0..����9do���|1���;,�{�[k ��x5zR�c�_��&�� -����U=@�RMq�0:���!(��NHON=~�6~uȶ�)E�@�:���D�w��f1sDYmӮ\�D CI[u5B����~T}E7�R<��a?T�9tm��e�ې��V#f*�"(V^L댇DK�j��m�4��Z��~҃:"g���`�}� ?.� ����[[�0
�x,��HI��Ox� ZW?x��W�/�y�uwWHhe���`�g?���	�&�P�f#�)X̏d-[�#���u�l��3�>�]\C[^}pn�w��K1�%v~�|Q�#d��¤vhխ�y���_�w�e�׫�k�{�������>��{�\� ����B�jP����%�=?��Va̿J;�!I�g�o�B`O^��`|��k� 5�ő�;�� �t�yKFN���r�^~FP�n�;�>夹�-���ϡ@�:�\���/h�ey�D_�n�TJS����a҇�9*2�������� �sm@��L"y�GO+�e7PJ�m*k��e���;���oO�9U(�������OS��^�'\v��N��Ȝń Ko��`���L0�|f�TT��g	vay����T��b�.g�����o�̘�����4�m�D���X�^g�+N��\4+����ת����?2� ��㣦[�����4{��`�^��>�S��>D�k��}r�e������%���3�vk��+�<�&���κ`�6<�4�ɸ*���D��e�\)D����N��(ýr9���ʦC��!�tQy�\jdJ&$q�r�v\���'(N?��9���^gj�HE�SE� �T����@Tֲ^���Z�w-�I��Ɖ�)1н��Y��+b�H�;�Ⱦۣl!Mi��Ε�HN����x�qCш��`����ZI�G/�#���]��[��T�4��T��;�ܳ���������1�*��	M��cUem��K�C��푊H�B/�T���lЄp	\��97[�R�%Ѳd!�XՀˡ<N.�F�b�ϭ���k!��p�7�V'��W1�b�n�T���>�)�fۧ.V�rԱ��_P{�X�kXY@8	1N��&��M㴔&�kb++/ ��m���F= �7k����-_}ą�G򍲳�.�{z����i�;Y^����P�j�Fh��2؇��?��*�:y.�藮=+t�~����R&�bk�D"NUB�͵b1w�j�u�x]��C6�()b����c�j,�R�n�V��F�pɽC��䟾v0L��i��6rFH��_����B��t���$����E&x������_#��N'\1�,,LA#��0 v�� x�^	8|��:���}�<���̱�C�]f���"�Ѧ�D���I��q�1��q��G���i������n�
88AE8��F7�B�3z��>�"e�/�$mV�}����ա�b��e[�y~?D��p�_��
���]$s���{��CtB��X�0�Ra�Q\�WC�-Е�=B{T�/2�*B���$����H�5G�.T��P	��硝d�	�.uz�|��ǌH��p�|�:˱s{q]p��N�K&xԃ��7%B��!��pZI���K�+O����g���@G�S]W���H�Ղ�eL�{[|K+�"����e�����;�d�౳;X�nI �9|��ۂ�$�0�q>�R���0|�����j��TF`�T��MQ+���0'ګ|%��Co�>CwFk���/q#v�������o���d�IFL�L�!�Du��~S�kg�����o��U�Ѡ����Q�:m�CY1�Kvƿ�קJ�M��vsNNOF�X��)�=^��E�:�wE��ѰMQeX!���J#��,�� tlg�Yd��h!:4sM����;��%�^i90׮�V�씓���{��&��"� `�R��O�=/�)����/Hl 2";�﷤?�����?�;�$QL��,U��	Q��A���T�E�����@;���g!�Ѧ7�-��#S�6�D�)q�X� H:=�ƮHg�F��V���6!H̖ rOY+q�@"m�bb��I�����P!�On>�ݏ�W.	i|nb:�$>�Ji'�#e��ǹ��AZ�>��@j��n����I�A~i.$�gT���&��V	�Xw^4�p�@L*���c�ȸ��$a;��ڶ�zĬB���f�<�Ua�w���Ÿ_��b��h�x�I��c'.4�t��k�w��[͉ë=����#x{��|O`ޔ�PT��u��K�2���&�������ͦ�h�c���*�J�9������j��T ��w_�Cm��8i��`��'W�
2��y��������`� q��g�|��5�Z�y =�i�1e( _�b��%���
y,�g�&?rh ��j4��P������)9g�R�g_;�\_ d����`�@d;�=��&.�P�qt<0ř������u�+�_��x�I߼��c�ǲҭ��x�� �c�_m��?��d������ؤ�4�H�Q
�XD�r��9i��O���T��ù\�娳)���w$�^ġ��W�N���	��F!�I�m����Y�%0u��|G���U����Q#���w�X����-S���M��������{�|�N���Oҩ�ɪ�i/���|�T�{٩<"ҋ�o#��>�����7}|���4��P0���X?��f�ח�\_ʹ��o�K�,��Ô�庎��+8an����B~וu.��`��g,!6G_��P�UT�T�2%$��_�/��	܉6�+遟�d��b��&��⭸ʟA�
��Y��a�M�B�~��$�YZ�Ϩ��nUv��}��<%�6[�Aǻ2� ���s�g�0N�:�ɠ+'�d��G���%�t���Y��2�\<Ke5���px%��ݞ!���>��y�3�
�-o�2')bY]�hl��~�)�^��F0C�iw�^��H��E�)B�FxN�<<�m1�)�Ųۺ䑅�~��m[��,�õ���b,�ϩ�:}Np;�����a*5c�AF���Ab�oɕ���	Uz0ȓ-��'5WcZ$��h�E��]W2"+)�N ��ګg�<���hL��{怓G��SA�1(�m#IS�(�"IE�v��]��pL39!���AVdW>�$�Y�=�Mc���00���(`0��L"�8�s��镉I�p0%|�Q�pj��{l]v������KƧ�>Dl�'�^�7������u�~���#.�Y�|Sg�n�}�Zk��s����j�[@U��w���'Zm��[ofdѓ�Mǯ��\O�)�fܭ�ss.21�񛵝Y9�-^7�=d`,�̸)�p*F�s�3WM- ��mF�ځ�TH���y�_I��˩��y�k	C^���#&�"�� ��  섍Yq_��(��M^�>Rȥхh"�Å!�|�q,iq�{0qĺq�T���W51t[���)�g��R� 4ˆ���+h+f�O8��d��G� �c֓�x1yoU�ࣉ����"�j�|�a���%z-'P0�`����[+�|�A�}5�*}�t�=m�n��~,���=Jn3`k�+�M� ������c��~���y�=m�cknM;f��!G���{�_�;+�8E�'�+�ƙ$�i3;��@��5k[�*W�'�����S��&�e>?��ڜa~��q�'���g*��>x�F��|��i����Ut��͇�y�P��\n��lb㾟jn�U�PY�.2#�G��D$�б�!I��|̼�Wp8I䟿AnVw���d�[?��a�$Ǧrl�W���Lf �'��ܳ�.V�KO7}����3[R�fl��M+���e,Pk�������/#��1��n87�%�h���|Cr�X�9���]Ö"�C���E�ٟ�Q�pp�d.����F$��`����T�+m3(�0q�0����Za�l�I�[ۿѲ�	'w���sUaF[e-Ƽ�~k$F�\(��A���4I�̵ֽ���3�G뚯��
���8�\AZ~�q��o&{Z��4Vf�d��h���p�=����y<C�ޤ�q��d�lsz��\8_r޽��K����=�ev�Q�&P��8Z�k���c&z�"?JRS���#܋�u���i��D���T�\��=vg�u;�B0��w%Ѵ0�%R�����.����3�}�q�)@�03Vv�I�_II�؇�C{������sG����́�e��pw�jl����U�`_��3�J�͸)�)����-�XO��=��V�����ej�켬ӵ* ko��I�f��wx����� @; �?��	�z6M`���"�X
f�3#����g���8
��������'iu�:��R��oކ�p�ȑ�aX��;<JƏ��~@����p ����.����$��F��P���T�c��i��i֠�M7+^��sJ%���X*V�3��_]f������������v#��O8����<6���e&���UM��+��G��+S3b��e�_�IA�"��=��(�n�KIV�˺���]r���ʁ���>
��%(Y�.�J1p�Ц/C-r�b��b�9���B��^u�h�	��>�	1�ﱩ�#���Rtzg.
���#�h���D�򪨂��=;���u��JY�<��1S[�$}qFiS;#U(�\��4$ܦ'V����9'/��>��eHKe?^�4�!��)^�%�Ǔ�5|��n#�䕂�lP)����p@����
����Vk��	F,���Ɓ�XG2�W~��Z ���hX}��,J0�W�7���� '���A�-��<��y6��G3�"�2���1|Z���1�K�}E����
�E��>��KN��6Q�D����!��G��m�����+���Et�ǧ�c�[ocP��oj@��{ș��(� ���o��}��;`�^b1J�5��F�a0�p_��I쾿���Bx'�	=��A����M�
>e����&y�h�?�k�>:�哫�V&E�ˏ��k{V���]o@�k��ZY���������
�9|�^����p��=��66L��]�A8�8�mxCN7OA�Rj�S��1��P�\g��:�(ďz8voE�b��|}6������5��F��2W+������ʄ�Od�1�S�kNf��6?�֒���\��<�Es�U��`5�v"�?�g��zg���쐫��!���$���o/�ҹ}��A��ġO�0�k�F^o�����"�V�5�7z��
�6�6);Z�bU��w����5��S�6Ob�Z=.��O�����\��m��;O�L�}��g�&l� 䬇}�̦���j��aq���j:q�����֣G�rj�\FA����z0 �]��v����n�J�ԏ��4[o�Kx��~�:&<`%$Fu1�KA�20�(��eD��D���@t#93U�����q�`n���X��fu��/~��9�4�`zO;RK���s�n��T�c�� d�2 Q'c�nӄ��1���Y�˰Wu���G������0��	�x��18�!�8���oR}�d�O��_����V��ij��(�į�x�Nݔ�́����A��T�H|*w<w5���`��0Yi�d���YF��a��6��;���0h%�_��3�~�%UDL�h�imsK\r��L6�v�D<g�"�6����ѺL��`{����2�p`8i��x<3Se��/<��zXu�J�GBޅ~T]�����(�,{��&����_JF[̙%h���@����5�t��+�ɿ����E~9$
 ���,����ڢ{e�LI*A��CXN�m1߆B�sԊ�vZ��P	8�,����8�J�(K�=�s�&��&����&�k��it����z>'�z+B��T	D4�yP�\��u�2V�*��45�4�7�틦�#X�3�Vʀ�)%��n��ɕ46N�/Sp5�䰮�I[�����!Ӎ�W����Y+�1����@��٣b˨�[�J;���3�X �StI�S_O�
\�q�3f�Ml�ZVu�_���F��Q�<ܻVǋV�2Y�~�������ǚ_j�[�(C!	P���+���@{e�䤇%�=Z�@#N�}�C~0��B�V��HЁA57����8&	���)�f`֚�� �)hır�b@50�-I$���Ռ���\�Z-�2wIr���_�Vt���5��g�A���5J���h򸠀�{��L�m�Ō6�p��B��^�nڨ�Nǣ�	}���6�ܖ�R��3��'�m=�q�Rv&�g�a�_���t���]�?܂&c�GqS ���1�.�K��y@',���v0�����W����v�RG�z�
�60h�O���ހȡ��ͭ��j�靀h�?��<�v�-��3J~s�2�@�ӕ��Њ�0.�(�߁%12��Nw"����v���?٣*���q��H���5ܜ��&�7
τ���|��)��D6i��P�]o���F�'�Q�0�X`*<wt$洔V��]$� �6���:0�eF	E} ���F��lJL�nN�Fqf==4�IGd>�:2����K,�r�p�Z,�������!��)���+��T���_���A��gtZ����z�Θ֨�A7�0�a<�������?~��7��+��SsD�]�w��.�wu�׷n:�����3#շ&�_��m��ۑ?��-��g^�B��󍘋ʹ�U7���IE�P�?G�Y¿�TW/>M�X����������ҿض
�zzi���䪆,͒ͬ�y+���Q�����üF2�� � ��KIX� ��;6�{�5�1��ᣁc��2�]t��U�8�j壧�F�C�E]Gq� �:x\�
Y�������J=�4��J

�C��D˄{�!F��F��Ӌ�*F�8:T]����b����/�b�ƽ�k���`5^�v!� �ɿ�	y{��y�:���&�8���:��P�dm�_�$��(��e�2M5� 7�b�/���[������9�8��4��4�@2r��|%���'��s�$z7�ŗ��y&��F���}�z�l{P����l0�q���%3&��T��x��爇:MD���uY������n��/��6z�Wh���GD�iۮ*�fP݀t�ՋA�7e&5q�w4]F��k�����,�𦭤�<z?,���PQc���| �>awܖ�I������i{�)*�GO�����0%����x���t;�N�_C�ڎay�d[�x��e�Y~���P�T�Nd�y�I~Ƞ;s
�OI�Q���Xre�?���l����vtyFs�;��su��e�Q�ܴ_���򥕨*+@�\���
r��#_E��|Ǵ�/�ҹ���A�fϟ]\_�Z�,ܮѧ�]1�N�'~�Wq�G�����bpMKB�(��Q_���C'��.K`B#|���z���n�Y�k�{�\�7Z��m�$2a�#aCd���r�2��XH����3c*�	h�̺v)����kK�YR0��eY|�zd�8(o�p��h��,m���MG	&-C��Д_�4�u�E�ڣxN�����x�? �.�TN]��K@/��+�ј�v��`���8c�-�{6���IkMC���+e/�Ъe먰�{Pﭲ�X	t�LqJr ��vH�yjq��	&튐�����w!��g�3
�a�v�A�8�-�aUl�Kh3��_� �m���Z{���\��	�ti�b-�r���T)׿߃�kC���Ǯ��k�4 ��8��/��t3�-@G19�i˕^�C7��J��\�a��ˇͺ��e �'>���[� �J7禟L���O���k�_���?�0o-+��&�����nH�#N�m)`6�v@qT&4��J��A�>�f�M+;��T�#�����
����o{�מ!����a�l}k,��=�x���w���$�_�K��z[�Q�����¦|U����>jZ�>I��bXO�[u�
�_#��	I	��Bd���S.[SB�\�3`^� 4�==g�8��`��_/ɇt�v� ���#�N$P�$�c�#{��A5ҕ�p%@Z�[N2�M�)v6���Fy�v=�Z�)t�v����ك����_v����p�0��{�ә�������r���w��땬J���������콀!����b�ز�À�/ t*,���0���ƹN&�}xJ�gP��^=>�+0�@ǀ���.i�8}�eTN�t��(�ؒ�r������$���޼� �(�����ZO�	��dkh�:.s��{T3a����1iO<�s�!x��˨!�x��jSIHV���wQs����+������ȑ�%� ���}���P:6fH\��	����o?V��`A��d��v��8�/l|1y�u����0mq*��ry�9�Va�;��C���!��p�����	ӱ�~
��\��+9tWI�z�R>�����#��Hf�]�a����fI߽>ˆ�Cq��FIN���+^ٛ�w8(Tli�
ū㻬��s�	X��/���E���ދ�+)�١U<,��1̅����9ej��O�T�RG��GGR��O� D/WD,0J�}N�%w.Ǎ��``Z�?Y��_�_rq^^�RT�1�6+|Dhq�&i6�u)�a?�u,ou�Z�?g�炤mH�<�;߰��f�JކA����Ӣ�qr�4h�&�������^V���o��a�X��!(��&Z�����,�
@)�87�_&�y��tϜ���W�XnC��37�.�Ԅ&66be0=�vu'P�2@Hu����<o����!�&�3fg�=�H{�Q��i=U*�^�Ё%�;�����D>3Y�}L�i��?T�[6�~u^���Ͳ�wm�5E鵼�|	�K:NpE[�ه���o0�g�$O��:<[�)/,�p�N�]�-Ăj- h�Q鐴����2���D�m@�ӵQH�.=	��z� f1���{E균�ʊ�Ø�1^�y�u��1}s�h�ו0"8￧��=���$�e���[�l�B�l�:W��������N.p�3� ���¬b���*[���Y��x�}e�1���;���m���s�N���b�֧��F�oo�ſ�6��w�,�]��a|�MFH��z�{��m����Ţ(z֫�:�\�*�i���@�Κ�����#�F�; �;O�崐ro`8.S�v4=\��~�m�p*�w�=2 	�a(�NT���ܠ_\��-��Ɲ�u�j|��}���}q:�폎 9�y������p%S��k�b#�Y������g]�OM���4a�u�C��B6�Q3�&�;�@��"5�r}w�Dhӄ
C�,�+��y�~�Ֆ n�T�-Q�3�����W��K#5#h��^������G��Tx����#Yh�Un��s��ͼo2�@�[��o����.��\���ƶ�����=o)O��[!�����g&+�t(:����TZ�;������Kh@F��B^��-<� �fȐ����tT����,���h*\�����JJ�W<o=�����5���(�Dn���~��=��j��2(��"B49��߃%���@�E��I٤W�/��^:������'ѻ���<!��@-F�u; �,L\�tE�&;�T=�]���<��h�65���|U�&�h�� ]Ap�
�r�-w�Y�4I����:v�q��z�LngS&(:�`f�I�$б"ٔ�DПZ\��43{�����N*���o�1��|]�ٸ�>���@���K�V���T c���7t��-4ʿ�`�������q�Je7�w-Y[�qܞ���Iga�����Nk{�:�4�3�*B����g����m����{�� 3�"ro�
�"*v��.WQ7��K�+"e�e$��/�I���aB )�e�H�����vQ�D�c!��c	&�d�oּ��~y�9.�q)`Ԛ�N*�2|��\�A�4�"���@�Na����g��W���b��a��8�^��.���gϖ�Љq>a�O���G�p�`�$��*��v��.����9N�5��h�R�mM]h|�r��S]�꒕%�(J���q���:�quIC����s^f��B�{/�y��Q@��9�s����Mp�G�\��gS�o�H�qs�ʦ)o��7S�C����o��?e�5�$R%�`���{s���Q0;����6��;ts$t{m���*$H�[n�Q�Mv��ˆ�=p'��Y���K0���%z�1���*�4��6#6��i��f�J��K��f���1S�$ ��d�$�-h8$���V �]�S��*]�o��M�����R �T�������t�b���Oi�.E���͜����f"�NZWD2���-��AՔ�%�W�p�d����%�^�~Z=v���5���a���U����ٝFn�&�t���Vr�xLUc�x'�l�����4�kX����}���(g�ę��`��2�;��	�&<x�W���/^���Y���Wh���4+�|hX��p1�8[�v;�Q����|k�7M�åt���֞svy�[��p�y�ULSXP�|~�RK�(�_q�J�H�zU��m������u����tT���V�m�T�������j�=���V9(�D4+<[�8��6�>��^�+�󅠊��wgL�k����PJ�Hԗo{)�H� �����yw�2�`����`2���7��ܒ�Jy�;�Ob�D���@��+�B�`�X�n�F�2\�<�q'��n��SZ�1B��NZǆ.L�}�`lDĕ����6�������y��I�TU�F��������F.���4x�-0ɷAny����j$�%_�'�8�:d��5���F�2iB��0����\�𺿲�,s��dG�{�`����?��G�&�[�-�[�L���a-�5
���c%@.D،y����2�=P�������(�!�r_�iZkU���U��������ͨQ�z�bZ�4CK�O~��r�:)�F��a4���X[��
 a0@��-�3�̸-��L��� 3K�����i$�~Z�g�������8J�W��� �� E�kT�Qr��d�I�c����PI�!���᣺�w��#�ƫ M*�e�ؘ�i��R��$�Z�P��m���N�G���l�TK��(�����8W�ku�Q�T)�3�LfF���G��	,j�����G��r_Df���������.��y���D�c�xP7�7�(�ef��r������`�\*y޿������ԿB�vޣ�م�XBH�/k���tYI����r���A�J$���vBz�0�،dE-���癖jϲ
��[�������.��N	m����˼T��D$�Xnc7\Oݯ�~���v�u}�"%�Ǉ����-*���>���b��`O�:�pSqZ���Y[=)���G���P[�:l]���{�l7S6���e�ۘ��JZ�>��������m��W�������>hdO�.��&�B��M;��� u���+�y-�>� q����s�����������͒|���@V3I�}5s�BOm�(��1�1J2�oQ�PP�jK5.E�����<�N�-�gr����!Ѽ-C:����Ȕ��|̤G��
�˱����Y��E�.`���y�`n+[���b�+��?0��*,wH+�,� �{�B<v^�	J�&��-b�}�B۝�fXؾl����X�4��E(N"�ayD*�O��P���π���BR��&�Η�EP�!5���XTWS:��d�Ն=�۾n[G��.!+�om�<��-�]��aы�TL���qT�x�;�?�����u���CV�N�H������D�xs�� �d�aL��.!;_�^��ٲw��u��#��3���ʥW���_J�% ��R�$R�w[~T0{^�>��ǁh����% ��)����8�תb��w��nL?�c�\�v��(��Nn11��1 ��=2�C��XF�1ȝ�}>�62��r#h�#3D�O�B��E.x)=x����U7���ot&"�4�>�:�i�~��0Ҭ����!��lT���w�����kЕGy�g��M��e����Yl:��Ck���:�� \ ��~;�1
�?���(��gJ�͔P�C�}�t�S\�b��gr���W�)�*d�V5�q���)�N�;w�)�>PӛG� �ZM��s�f�&�dڎ�o��)�M\��K��aaf���*����^1�z����qNU���_����l �U_��I��dt��
(3@k��k�
CL�a�s����x�I$�s�����an��c��k�X"qlX��X�x�8hd���$�П_.w���Jv���v� ��6�j��R]�-�f��*[��p�m]&�>�
��*e�����A�(������-|�4�I����w[ĺ�����S��P�<@�+<%n�GTJӑ��d˅5[5�pN]O�4q�Oڅ�W�Ů�i�A�|`aL��B-�`m�o�Lj[v���7n~�Y�Z�����5���I}�Q*�d�c.�}
-��x�;0�F��
��)�	hO��8��6��rc%Pi�?衊��&Y�/������G�ļ#x�_�ȚJ�ᦳ+Cp�|K�	����eG�7��{[{�e��0-� \v3���Hs��|���+�E `B\��SE�c��T۱=��ĊS)�:p�y:��5�1y�Fə�s�
���'ʀ�q F��O�Ϝ3]\ܼpi%*#��[���`�5��'$�p����6��M	���.��v�,�>F�J��c�%�t��RLc.l1��A�R�e�N#^�d����jY}s��COb<�J{�����D��WĪ1c���#���� �3��J�Ԙ����_A��e���4�j��pl�.h��0J6����D��J=|l~��.r��~�#�Ɂ>TG��J����+^
����Q�7��o�e|�$i���[�*��M#N� ;��m��|��A�9|q�n�%���f �qy��FAzI��9��.�j]��	�����(�*�k&-1-�Xz&
�1r4�y�`�ILt{�0�w�,��o��M	]	������W��a!�
�]���.Y�MM�[���1��?�~�r��"Po��|]����h؋�D@�a9�ˢ�L/����W~IEWW.�ٕ'2��|��/��_q��g�J�@d
І������;17���4�9 ��������xQ'�	V�26��i7�z��B����J���4�k��ؘ<k�W��,����ڗ��D_aS� ��ʕ���?�J1w#	�'R ����O�6c҈�΂}�MH�Rg�&��jW��}�Lq���~U`F~���I����'m<�u��W>r��@�W*)On��Z�Q��ϖ ,j-��uv�� R�*��ж��Ԕ��P�� ��0{/nA�
ɢ�k� ��>D�)�[.%�Ӌ�*/�k�q�/"����2�X��{33�w?�!-�zI���K�5�V�s;�!��4�wR"I��H0P���:z�fX���I���@�b��a_1��p�B�����Ԛ�`�]@�<M�pz��q������'��
�Q=,�n��d�� {4���h0��56��P���xį_�VN'�y�º�V��}��w�� ;ǆ^_��>p|��uM߁"f����a��%|��ʼG���\�e[��&�d�8l�Q����e���u����rmSͦ����_>^�	��!�T�𲣻�64���ׂ�Y#LQṣyZq�w#j�@���H�L�]d�Y�S��>8lܟ)��BZct���>�:4ݼ4��m���5�8B4�)�ɍ�\��L��p����mƟ��h^�E֔�B�M"�bG2�C?~��Q��cBݓ��U�A���?�Z�^xzr,U��-�ɕ�� ��4X�c����g�wmc���`S+��G3�&ۭ�A�)�~����,!�	,�¹Rp1������o���Q���*=N�~��	�=�o3&tx$��+����][ �V~�層�f�	wk1$>ZF��;�3U���m��U�u
�>q)!�{�d�:������d�s��(J1=�_8w�~)�XU�-��T��Q'f<�K���[�1x�wѷi��С��Ā���W�����%���WR���w�S_��%�-��ne���y����R�Rq���J͓Qͪ��u��fM���܎��Pq�!԰B;����K�����ȭ��c����]&���/~L|1m������z���w�)���r�/�+�i~�5V�z8���BX�^���n���$�q�ŜRGk�Q+�_.��(��BǕi��=xyC$Lh
�A8�8;\\���cSe��%:�����`#�wRh�|��H���2X�,����-�=V���UOo���^��&��a,o%�G+xI�9��$*��a���:|U$�Z�}).���p� �r�V�&�1��Qլ��[� ��k��rv,����'c�X==XyB��/�ޞ�K��[Q�L9�O��F��E;( @{[�k����~�E~IL��GT5�+gʠ�E�\nxN���l�SSX["�mh���x����\;���5����w?|�����c�\}�s��`x0�|j��X�]������(r���Ub~� �V;��˵���`��~F�9n��E{�Ba����}���!������U�	��\��[ �R�-��ʹg�
��] SךXŐ����K������=�C��U�'X��̿�(X�s�J�|���<|[�~��;������9����A�&җۢ#N�J�%�ʄ&��Uڂ(1��uԄ�#?k�W!d�TS�Pj�0�ꢁw����������,x�H}�[������+�� �{����W�����Y�Cj�_>��ɱޟ*��Q�3��DXT�b�hn�����ny}��&i�����'D��o �D�&��÷$c���Uu&�K2#�eҖ�3��6�ѯT��yl>L9N=c8����s�B+#���T뻡���.���Pc�#�sT��0g,���S<e�����ʇ��9��W:�x�ǫ!nϣ�Ŧ.O4��B�
cKA����b�aP!����nhY/���p@�ņ�V��$����>X�y_�e)�'P����6��1��S��
r#�=5��*��J����ķ��{��U��K��N��-_S�x񪅨�='
���3rC���{�~l ��?M`q+<^O��A���+����Ճ�����Z�0,)�����s~���9��Th�uV����Ʋ����?�?kXM��p6�a�.�i;1�t��)�_��U�[�����;��(|ir���G�K��r5��_�ם��%��U����q���������P�@fZ��mwTN��,�ǻ�*hv<ӎ��~b��ט�A��.���!�"LW>�m���-��B�.9:��A�Z/� gҪ��ͫ�q�* �"H��ŵ�fb��(��h��<S�9`wz~�V��ɩ�T_U�N��y�ä⸶�F�1�����`�ZA^��V�f�O��6.�H��b~�߅���/ir&E)
ق;��i!��"،���&�+ٰ���I%AT���`������q{0�b���������N '�ݩ3 �GYX����Ā(Qd�?/��.�w�k��T����\���`�3S�KG�f��,�уD��+�P�?n ����3|S.���8Y/q��6�ݣ%w!��ꯁJh��huHM�U,���Z�?Dg�;C�>���٬��Tö4�'�7;���H�9��3����nw3H*�$�XY{)0E�����ѬR��/�Ά�(��>�&�v�P�-2`� �����&�����<��!��lD��Ҝ�a�+�����{4����i��`��V(���UWҀ�����Aa~ ��Ոh�.���ڿ�(�P"�8��㒼��vIk.���pAƂ���̑@�.�&�H�9	����.#3y{�[D��k%'�.��(�� g�q{DsO�}w���̱V�%���ҵo���n������+ߟ���R����Q���C��P����#m::~�� S������V_�E8�!ـG\~�qF��w,�j#dnSԅ�f��6�}:�L|��|%�j�$�� �s��+�b��)�D��ucm_n��^zZ4�֞�p ��� ��[���@ߔ���� ��Đw0}�����ѧ��2�˪A�+h{gؖ��S\�0�qOH�o���gh��ƪ`�7���P���C���Lf��ء�����$k�I�N�	�y�8�9en�����g`��
;T0�� �����3��+�^�ȵ~��P}��wEsm���
��T��X?�є�8�Q.2�&��H��Z��Z߻"1[�J>�9~^�$?T���򔘲�Z�%�E_�ٷq�n�C���w��Mt�lu�%��L�AJι��	�x�e�1dF�\�PϮ�c�v�V_�S�b��{�Cs�뮉n�q��^3$9ϑ&�Z�1��*{n-�q�u��x��8���A�9|�����������A��-���#B%��|��7_����˫�9^���˦��#3����tAy����T��tq�h��㬐Ů�b���\0!�W!/X�$;��/� �9�.�죹����6��8i&k �7���E��^ԫ0ꂒ2d��
�s��́V��iCS3��)Xܵ��f�����	L�^�&U��:�m%�Jc����K��F�����5���-v�J������qw&��D�K�ER�����K��i�0)7T����^�6~�lO��R��A�	Fh��\B���a5"�o�ȝ�,������
q!�E,����P*��'�QmpV���wo����;����E�ҥJU_Yw����i`��sA���h�Y��!�4�]7(R]�.̣i�pX���7=7���	K�BA�@s��f�����}�1�Ǣȣ��+Ro��}�O��:�i�~�ƝC��$��0�����X�u~E+��u�I2bۨ�48��(G�8)���D4�R�K�㍴�����R�藭 䴐Մ����]UNa�xr_aÝ���4t�֔J�,�!���^3��U�z'A� ��ryAK1� ��}����ԯ����Vo	��X�!j&	^:�v)cB������'���[���,b�BpPc�o�^��ǜ�����+�`A��ptMz�!".�m�G��]��i� 9���25�ғ� �y�0	3����o�0҃�c8����ݷ9|��v�a�w�*|b��^l�n�鑏q�_�.����»V[W��C9�B<�
r�l����o:w�-�t�}�����R0I�]Fvfk2��hrw�z��$�8J���ѬE�d���u�ү˷%�QK=hH�Ply�?���v�,Α�/{�ς�gy!�j���U�K�^p�m�x�М~͟[zǾ�Q@�g�M�Is�|� OA�%��/�tG7��c��߿�M�d���_EL���٦�:j�x��5N�G1k�d	�h�G&kV9Mo��F)D�P��1,���\�dy�9߃f�lP���é��lZp��T}D/)o���Kߋ�N{q�����@h.2ZE �1 ���Ri�8�!���TPue]�^R�����h9�}��zʯ���kj�
v��,��뽐�w^"��1S����id�Σ�C�@���I:�����T� P����w�g��#��ߢƇ�D����.��L �*PNK�'�Xsq�5���g��[\M�u���C������ C�HЃ ��6�N{�ۮӊ@�v:�ʰ���>k���!K6�AI���AS�=�?�d�#/�
��j)`C��Ck`��aCi"�K�S'�F�[O�0��5 O�ڬ���Ǭ�:�F]�S��4]��j0GB�v�F�7O�_�Q��?/�H"v���*��gt��)U[O�Ҍ���Q"�����s��NJ���#�u��˛xӇy2<�d�p:5�oec �J��>��7:���ģzlhݎ�nտ��7�[�W<�s�d��8��C�����o�e$AMN�4Lh���פ�^��W�}�HQ��a��Un���D����@�U�����ZyÇ5a0��?���]�
��PP/mk&|�e�>���B��w��s���j4�;�*�?Q)��V-�i���qt�;�Ŕ��C^�<�[�I܇"��.=lb�FSP�,���9�
���}�f"�tI�AH�:��6�:�}�����7o}�p�Un���y%�ZK��kcq�mAIT�I���t������ �}��4�=�;������]o�Fք��r�n4�2= T�a>�,��u5c����*��DW��kÊE��QI�����5��@�%�t&z��'(�W�w�2�`0u�>'_�q��Et� ��&;�o�Cꃜ�$�:�E�'�/N��9D_�u��u���lE�i��;���Nţȧ��J�o�?'	�ΟՐpi�_k�2ֲ�_e��jk�d��h�Ɋ{W���w����c.���L#�wX��P��x�[����_���y�T��k�
V�E�ܻ�(2W�j^/H�L�h  ���p�~��]%n<�qǒnM�G�����b|{%��7���XJev�~:��e/|8�+��7U34��������^�k��jK���i�۱o'`ȅ|J`��/_�~aWCt��ߝ� 		/�|S�����#î�{eS`�	�� <Ì����r��Pw����m[���-d�����	��q�"�q?��r<��7��
Z'vzM?
._j��ɯ:�Y;H���N\�M�u�abo�&iר�!.bE ��:	j�f]��@�j���E]��bZ0
S�GS�%y���~�S���a�ؠ-�>5��)}#p��g��+�����Nr&�q�	�x#�фz��{�=�ජ���ziX-)�~"$�,a��qK���YL���x�;v�bgX�-�i'��i~��Y�'+����L�s����8�GeK�L�LXB�s:�+�`:�I�d��+��������Bm�p��OA\��t��|���8�m�W�uu�W0D�S]	L��2�U��3### �Y������]���ӳS������V��͡wer��@�o���6�D�?�$�l���R��vi���8"v��+�\N�s�;&I�xj��s�����G�{U�l�̠���a�����MB�ܑ,Zv�'�]@��}�z"� �,�����f5�"Nc3��!C#��A½ ��'�iF&k��F�we��M�pl�+��ME*�^Nf�D�Jľ��Pu�3�qɄoe���&��Vb<��Z:�(ߐ�0��k�%&̱�!�D�?� ��hp>�W�)wQ�Qm��9��$c���3���Al�.�M�MDzÑ����|��^_~ ���#��'�S�ĨS��S!�Gw�qVI������$Z-�zG0�d�c�僃�3��b�����R��i͖������I��k�h���8���p�򋀤HT�<��IH�&{�]�b���C�.�T^�-�'
��E�bz��@(������n#�;�!a��5M��e�69�ZV�?�]'k�@3�M��Ug*1,i2���f�~C�e�Z��,`
ν&�$��P��=�z����&�Nj�0��:�P��T�n��I㮕����7�nE�<H���-�ʢ���*�Hy;�t���Y�g5�1�̟ۑ�;��c���e�ho���F�Ck���|�B�[<��0	����RA��j��Ȟ�);��(ri�vB؉\�6�Ĺ�|Z�bTKұ4���K��~��܊�;���yR� \�''rH)Kt�1
_^�ȥ-MU��Z+���n��Ê*�a9�}~��Ē�4�n٨�&�t�����#<0�SׅUHgF<�dS����u���&�+ǈ޷M�5G7:/ĝ�p��/ou��رt=ٷ�rc��k���eӨ���L�cך�`�;���C���	�|��w��cH��0ю�7�*��ba?s�2^";u��ohS�p���?m��ZE#&��ɧ��M)-���Cb��,w�ET��#(n�߫��=�i�4#]dG�^��\�i�\����$��倣rO��W�e�9 �#�6��4L�P�tU��Nt�-�����D�UH�·��5ɦ��!t�l������%Sk>F��k��h"t�U��BΥ�'��;8
���h3��^�c�;~v�Q��<��,�9)[��?D/��KN�"��i?�]l �F̼R_� ��&
�����uz����gX�G�3��mz���^��.�ɥS��r�0��lY�j��X�9�� )�6)|>Ijx�g:۶�d�u�E+=0����Ϊ�˭���Џ��K��#W��D{��&�Џ~g���P�/��x\�8WR���Z(J��i�S?�N/	��bm��-nW<���x��n`�����_?_�Q���6�v*��IK��AB��
�����y�!e16�$����i*f�EH�����i��ـ�Ӱ���42ݫ��-'����8�y����?3��	���X��R�H��i9�9�B�|�P��?��Lc�zj8d��G�۷MǬ��J�N{�kWtm؞@�(�ȺaM#�Mt�,������j�$%2�,��fV��s���wɕ���m܀閱�G0B6�:�
�V��� ��p!��U�S�J�<�[���nÊDm2y�����,Kf���%\�r�tO2����<�S������� t�\X�&a��ڡ�͝�e<�z��j���gX0��z5�'6Ͻ���\G�p5��X��oz6@��TѣqS�Z�R�����Ʃ6�7ܸ����5���mv>�NO˜T�?.ٴ�#�S���}������Ϛ�;vX��#U,��ۭ2��
Ι��[dэ�[������	���A���_$h�CwZ��fr�T��ȃ��s7��G�6�t�N�>��@:r���v�em�ҹ>^AĐ�[P
�K�/ݮG��~�9�Rü��L�h�n�X�:�m��S��S���f$�4+���+r���,waϸx����t���)�bhLZ�����|Ah�0� �1��/���)Е�.��SVRj�)���4�K�Uߐ�|�Jt_Y�9MKB�	
1]�B���s�ȢJ:U����C��ڨ��W��N֑�T�"�yVw��Ζ�5K�ޡj��BMS���6:��!��+�t����x�V"�w5ř�	6�~N���8Ao.��H���y�azڵr�R�"֠��oAx��!�m�I����-w�=��(
k�)td�Z����l�����!�-#�!�3�`K�����.1F�Q�ݿl5D�)?�ou<�bj�N�����S�u�`����Luaj�w���C�#�ZT@�ɁK;,�b�V �L�҂m��<�z�c���.blߴ잎V�U���ET�"1tl��39T�&R��$�B�?����G�I�I�q�]����E?6Y������N���"T��s�y�&�#�∔ p|�Gց!v&Q��?���k�{����M$�Ab��).o�q^@�a)����I�=�)��x��?�����F8�7�*�.|�����=���`Wb��8?!�s��*�K��a(��)rw�r.ѷI�wG[�^)�X⯅���s	�F�h��G�j9L�sm�o�ݐ;�t�^X���c�ٍ��wa]0zb���=�-p;*����H�dxc�y�e��l3���4�&�a��Gg�x�l,)��9�E���2��W�Rs��R��xq?౐
Dy3�*P�x�	ٞ��EO�Y����C���0D�[|�������Ar����1N#�qw��&
+lH����F�l��U&A$�k]л��(��ܜ���,�}f*�Պ�ٚ�ޱ�9�h~�YKZ��	�/����K�x�0͢}7��ovu,���t�%��E�l�=ԙ��돾=ɌwD�tIȦ��-Q)�e7���&�:�c1Ϸun|&G������e�\���o�&�`$�i����底H��k�Ha �]1'وh�·6d��2��]v��	r�"=�@np�FY������"�$lR,%�p_�Z�;m�K�8�|���*RJ��Q:��)��_ݺ����@��wJ�N���;r��_�&h����9�����c�6Q"�͋U�+�(�)�%�z������
�gP�i�;ys�HKmk���8�DD�;�	P�n��#�t�t��ڸr�e��9cF&k(JZk���T$-��Φ��f�<L4���q<yn�g�����N���}w��҃vS�����"JG�`��h���"�&�0��q����G�L���I� TLP̈w��4��� >�U�́�ٻ9�����T��tw�.�Q�\��0�����$��Q��_�$�����|����0��R�oQ·�lڣU
����P HX� �y
'�S	] th�˚Nf<��5�2b|���^Ah�y�!�"�0�+��E��O�X3^����|��;���	Ĕ���9��P�=e@�"h�b]&�������z��kk�\Q�b��~l�s��c��WTR��Ȓ=󁫀���㩪�e�V�|�F=E!�a�oM�/i�a��q%��d���3�@z׀�����ƥxWe	��u�_�����nޱ��0�[��l��L��^<r�DR�g��.��\~=�Q�TQa5�U��*A��u�_�_b�uV e�>���JP*���1�:�����ů���h�0���o'l�F7bҸ��VD���\�1w=$1n��2X�:����is���	�Dg�����	Ew�٬�t-�>n�CI=X����,쌫:�e�1�ޭg{.���`'��+tY�B1�{���=��z����|�_RB�����C�ms{�cܰc�~�m:/�oz�w?�;h��;h�2��|��bO�yb�'�����A�tf5�ݫ�<Ϯ9��3%��ȕo�D�"���T�i�[�����:��s��D�s�f!��vN�zX4� F�z�����T��:�^����s��mQr��{���揽�w����k}-��F�6Y�d�-^N�����]�C�`�Fܥ�"$ȗ_e)4E) _��B׸~#���T�ِ�9z{T�i�O���d�懶w�}y�LSj7��	��'���P�س���l�6�5$��X�xܨ�h���"�8G�Y��uV�t���&�ի�5�aN���a��G��E�'���8��6ɯ�H��iØ�V��t��@�k��0����%?m�0���y��ñ֧�Y@���01'������W�ׅ00G֣�>����N��@��[���U��Xp�@l�����e�L�<�׊9/��!�)P�qw��{X�r��x���k<�l�)�	z�R.R�U	l�T`�\����K���k� �f��5����l����jP.��D;=��?����i�$w�^��s�./�l�"!%��$%��.yVU�@��/��Ћ��0�OG�Q�=�3y�ϿD04BM(La�8��A�>��6g��m_�H����H�SM�==��D�a�TBC���m�r��MU�p��J�'���^]�oHx�@R�# u��p�=�����D�v���Y �<�e�h;p�!2.<�&K���	FH��k6���o���5�ݸ��uWFs"H��W�.��S;��N)o�p������	�e�(��ӔB��g�o�8E���;3�@m�9���H�; =;����N>G�d4*��]>m��7����V2�!V�G+�?����3Ս�u:�h�@3�A*�Hc��T"��c�Ւ�`+&����s����TZ`8U����/y�Q��{dwi���( ^��T��T�&\JB�J|�P�	�1�̂�8ћ�;_�r��	�CP�ھ*�kN=��Ӹ �� �yj���a'��)�s��@�gX��z��g�!���.�m^���kR�w�m����`1�F�G�����܋����^�LY�L
�C�	�1G,�-.��0�\	���;���_tYz�5e�o����!��R?'�����~��7[��,�%J�S�ü���0�"n�pi?�E�o��tk��s�*����E���V�#�蛟U���5�w5���&?Ѱ�p���3 weZ���;چ���D!\X��<|ZU�|�5l�\������L�_`EbzG�b�i��N&f�X���w�ɀ��B՝����72���<�-+f�r'D��4FRr��}�
�����>"=\���)�a��N_��ت�'x[�L!�RboL�{O����ÿ��@��K/��NX�Fd�=���@�8��5c�D�Y�ɥt��g�=`�QgV�F͍���EP+IQ��(6��vPY3�MA�;�(���[�vb�� .�U7j�p�;�B���������5�oh����LZ�#��@RXh���)h1��;�Z7�6B��]�@�5�:Z*��ζ��>���~�oҌ$'7��?���K���Rw�s�hf�ZdN�j�X��Y�ިk?�ē��rH�����n�Q�Be�dʕ�� ��(�i�+�S�x��5��
�Gi%�ꄔ����M"���Wk�]��d���T�VskP�ǔ�Þ��u\�"�YHT�%ZC�Ɔc�y�$t57����B�yՕT������S߅Ƣ���s�i��A���M�݀R{�xl��Rb��t�ʪ��(�a�f�R��(y�5�HM����M�oL�[�RBoG84s�?��<��f�,�����7;*25���ʞޚ�q��rf��OQ�dχ�]�����E��9&M�8����ѻrL�V>ݬgu}4v3��6)�b����[(;ڱ����2�x.<�I��Qk�9�A.��jP1J���jf�4�̡��$Q6Nm�uP
��$[&CF
G[J�z��#�P��M�rfl.��-�B.dT�����ޠ�sE!+�r��z����3�h|� tu ����r�WT2��R?����B��]X{avm͵�E���EC�"�a��$�D�u�����/'>��'�� �����t�yo�J�zw�Q�G��\�s3�wce��eR��@�J�8������� �q}������ehs
��۸������7{�}lg]K�.qT6�ZবQo�|;ߨo{T9�
|�f� u�#�1�9� z~嘳�F�l��L�\;e�K��`~W���"!Y8\�eN�s�o'��n�9�{�FTH4��%s����d)�83C���CP�/���L�rm��n���~� �_Kw�C,ذ��?��PK��;J4k1�:M����=Ax���4C�M#�5@­�����8����4�U�8�-/���|�қ�Ջ��y���,�!��Kz�K���n��|��ґn*��}����{YZX��R���2΅cAǮ��Z�'�����Z�'I8R#�D9��+�.�܊L�~���Κ9��д�,x	1 4���{�c� �������J����iC�E��u���O�:L���1�p?C���Ge}B�:t�n��"J��V��K�@��Rq*� ��kK�|�w;,T�j���@���.���%�����>i�e��|k�i�`�"��ƞlT��4Y�>������`[�G�	��w�Ui��C��ö#^g��B�q�1���<�މ��g�}���in�v�0D�������{��E/��y/�>�^�`S��]��=�@�檓.�v�܃23��y��,�^������ژ.��zo���m"�eC������8`�;A!Z�t�c��|��E�Fp������1p������s�'�͎a�p�^���dM�>�"�wF,���-ɗ��.���_��3^t5�g����NfL�U�,ӊ���*H�.���2;�x���WזG֎8��C����nQ?��?�+������#�f@ezO�SI#��=�Q1#X�X�i㳵$�Cy~S��8���j�zlnQ�����]%O���_�~��W¯����y������ؓB��H����r~����_���?ڎ�11O�9��?�9?�k�X$��~�S��ԁ��M}T� �d��Od�{����(���)�ʝ���`���0�}Ѣh�X]�<u�|�>&Z?o�2QR��1T��>$�x�i��m�|��� H���]*$��P��m3����V�)��)ؕ�R9A�!���S�
0sS�t^n�ֶ��"%�v1��S�b���5cXG8FX̖�b�@��Ұ��ֆz���Wr�$�f��~^�����vʨZ;	^_�����,�2�Ô%��_�y��֫�%z���s�&jܼ�Nw�h"Ֆ�Sگ��Y�kk΅<Nǉ��
UrW�8�銱A&	���H�{�q�;����5���]EX��|ЧSk���Ec�����|fg��Wް� ��W��eY��;��o0(��y�RP��/���t�$��ᇐrR�쥃�R��z�uk�C�����v<?��*�-r��o$p���	�#�5�����S/\�L[��� ���5U�ʿ��� ,�Ƶ�2[D7�NqOƕ��v�8�lx]C�8?P��f��KS%X.u�	v�.~��&5-�y�ӞC�C�>�wQ2D���u��&��/H~�40[���P�^H��_lg��n�����ň�j{^�U�+}�Gڹ!!t���4F�#�]K3IBe�ml�6a�n��v*�ЂM���q�� '{�JS��'/�}H�f�ſC|��vcY�.��"j�&X�^4ԁ;Ʒ�
��Krﾞ(�oȝ����<���������[3�Ξ39��6rY���닷LP+|VJ���r�T'뷑�Ϫsm��������P�����=`M] A�d��]((�}�b�xg���(+J.t�:"ԯie���F�)���h��E����7�_��=>��"�8�������o#J�%��6!Q�j�~*��o��&��&Ea��,\(3�;!n����>=�̇:�0h�	Y�� nj�b�_Ca<�@L}��˚�ش��$�Y(�h$�}r���}"Ul����=����#Қ����9y+������[s��&�Z>��A�ƫ|�d����%��Òpo8���i���n<��v�����O+OcҎ���z�bLM>d���TSL��&�Cߓ�b�R��i؍��J�r�U�@���Փ�sU���X�) �����.o]#_~{ڎ�ӱ�ۄ��M���֬�]b�`&�5��8β���CU0�ԱR�k��o7#�x
r)� m�[�5 >G1�����C�R(�ȲP'�V�yM�)1�������4�ꩰ7 �����	;���B���N<�6�)�~7D�8T{Z�7ϲL�g�e�m�&���5ѭ^�rHD|�~Qҕ�ٕ�ȯ�  Kn1�#��}�Nƒ���]
7��LxJ�S=��𧉻B�HLW�w"�������ۮ�>,OҥVE�f Y�{=������:f�a�4F7J;'��߉��֠��2�"��8DP�؀��9��}7m���h�'��%Eo�.��d���z_48V$�n��寀�6�Mv��9	�k.-��P�:b�2�O���	qo�&W.x7�'fZF�'��d�]r�5�: ]Gl@�%��n��m;��"T0.�kR��Q��?������h�)<��-�3ӻ�`��D�:�
f`(�*��E5��t+(�p�)�=��0�`o�,��D�ҧ�}|��$ʉ�u��h*~pzM�C.��\�ܝ�,(�����������U��$l�P��B�&MG4���;��P�2��l ����G����^���`$�I�W�6��/gU�!B�~�D����}N��_�a���Ri�{�$���{2�w�j˟d�r!)$_ٰ ϥv�uiO��):��� a�դ��d��j� =~�૛J��HN���t<'e��_��S'7���$yG+����b�7t�Uq��06�[�=N��0a���`��S�I�S��f���
}�LX=�v��Ԍ�We�y��շ���&����E��S8� *Ajĺ��X0jDm���.�-���vRLNA�h��icx���&to�.lg϶E���,�,����nw����_��/�G�sF�b$�J�@�����]B���N�T����f�nz��x��1!�noo�8��fq��-Y6H���A���V,@���`<�2������'�!F9�ǩ:ھ/�{��3yj��G6O���Z��w�?I�W��`��A�K��.x3E� \+�Q}�耆��W���"���@�@���ۅ��v�~A��+>���LV�5��d���B���d��gs'��Y6(�n�y������8�$�M�sܠ)!'�KݱKiշz*�3�)Yb�(>�� D]�����;ZQo�[=
-v�Ư����*Oq ��/��>�6`���A[>A�Q�ܽt���߱�g�ܱ�+,�ɳ��Z��60�_���蜸�)�l���</�����Hx���v�g�X�+�]�5U�S�̒G���V��stx3�����ELdV���R��<�#;���0����o�%���2)��xsgLE��Do�]ʕ+G9��I|�N�Y�-V��ȮvU�\~�M�2��u��[gĪ�gCT��aŨmz�;�0u��<K��/Ⳁ�x�f��vS��s'
�<��dJ��WE�;���S��%��-\ˇ�^��h��]�oΝ=a��T7������ܥG�G�DG���J���k�A����47�-��}�����;�ㆸy*�Ӗ���{��HKL��F��
��ϖk����
2(�~6�<���M�}�AE*2�A�Y��S����~KY�m��tR�D�+���9�u+��Cj�M��n�N ٸ�h�?��fC^���r��Q�[�u����	�%�"} ���ʺ�F��1�[��7���E�1wǄ9�9ZQ�������!�U����	R��[�L
�+S(V�r�sF���t����6'���$k$����G���v,���L��.=����V@���*�m�Ƈ��G"��Z�S|���l�[�Yt���O��?	����.�P�]o��r8L�*��w��H,�1���������M�Ʌ{���Ct��Z�]�`���H��H��?<�����S�D8����F՝rR�AlL���=���.;�9^����͎�?�s��o�VC����>O�@�M��~M����ͮ�f����~s�������JJ7���9+C��	�T�%���#O������X�����F��r��d!��0Ԑ˼&Ш=;\��B��ߟ"HZ��3d�)ȇM�#���dG��F��R���Г�"uc$#K>�o]+���R4�'�غ�̦<�*���?��<u�Z*�q���:0m+���)_��=,��ymT�F�XБ��lnm嵫����n0M^�%b�<��^�V�����弦s��&��}�?jjKP-���9Oƅ�$4⥵��o+����֍ҀN@�1�(-���S���J�Ŵ�Wx�2��6�\-Rξ�w�����!��u�2�Ǡʯ��Ā�ಷ�n+�>N��3�v�A���"���V����@� ����	~�D*���ېZAű���ZE��>4���2�o(��tD}/��D*(���D�6�#�2Ʊ��O�������7�D�Z۷ޑ��w��Я7�h߂�dw��G<�����#\Ǳޝo<G��֥v�A���RqC�:�ݸ�����TE���$68�%m!C��[Ǥ�]d�K��8�n�o?�$�)w�y�asQ���ӫ`�myż�.E���Շ��g�@]�Sc��g`�Y�m;��������Xݬ�-�/���q����L�>ħ��-3�lgzi����"rH:l��.{g� %d!o�p��M^%$��&��`7
��̤�[LŰ�eI��C��z���%����M^�4��݀CD��笪��Y�`򽨰6���������c��6^�v���i��˚[��z�?;o��LD7qv�P?Hy�ޞla��*9�y����䪮��TG��l��E?�u�q8�7UJ��v��C�½�/Ѿ�)Ѓs�U�O�<�ޢo�s�nQ8DoY櫺� t3.�R��s�Ń�j� u_�j��%��|�q�?�WC�|m0�b�紮Zq��id�/\�$���Op2@;n�§�d?2n)h���u/IEo�S��#1��'oZ��/"���HUb�O�R-�|�=Kd�H�U	���V2,�+Byar�JH�S��OX"��펮�n��.�*�A���K<˕5̵nht�ڒJ@�
�B�r�$Y$����'��~�,]&fbH�	�Po���gŤo�m>������������WD�O��fi\����')���ˠ/�i>Ge�7îf�JJz�+��$X�q;��.�Ɯ���,�����z�ȿOg�:�N����G �����x-��@\���ҥ����<��}��?�(cc���h�	`�0W�$*� T�0M��u��3�f�Lߗ�߫��D��_%�����Ɖ`E��?�+i��p��˕@銪1;��_�U�ޜT�3�sׁL�s}���Cʧ��%��?N|k�>������O�𦦜�M|!�c��_Q;����!�v�[�����l�plq%��Oq�-wR�d)���C)U|��sϽf��LF���9|��|�����UF�Y�Qߦt�V�������������'�c��8M��YQ��m~����?�2��]K��9���3k�"��E����/�D��-�%	�M�	�ÂŶ#	��}8�{ s=�˄@r��E�ۈJh'F��ߘEWE*_���'�"ry�{L�|�}�sm�Tﾚ�܈�(��\�ѯj����Wg
T��p���Q�e�ay�Ն���eF�Y��$�gJ_�P�iY/=�/�E� ������y����v��6�PRze`y1Q=:%��8�L��{�X�Neϟ�Y�j��_�����Q��x��>�ӡg�y��#=���l��N�R�A���͑U�Ym��'֨�m�R�;D7�6<_�3��k��=Z�52������������Z��b��Oǃt�?� 9�Y��EŅd������{�ܛ[��𣓂� X���Ö�T�T��k8���E�/�	���>Ns���`gv���Lԇ�	�cΚ�F���Gw��g@j���"�Ϲ?��Q�z#���N��H�@���%�Ak7�qϑk�庍6����p�-*v���o=�}t�[��ltjK<aT���"�ް�&m��lA�D�U��bA���N4,e�U=Q?%�AL�-�UY����M#��x��j�5��-�V�Zl����~w��p/�@�̌������\���'$�h5[}^Ah.2������^<��<����N0\
��^xjm�5��R>�!��;�)��@���9��t鰍�D,m3yQ��Lo�T�H��;�wu�ӯg�|��� j�.y�)�k$�����=�
X��H`&瑥�������OFuߣ�3ڞC����c{P4���QB�	x�@�X���IEiG��0Jmst^f�v�����1�S2O�Xgu��t=Gb)��3��0=�=b�iVB��(�U"�|Oz�v�2��P���(P
��Y+N
�λ�Fji��Ly~g�k4DC�k����Iq;�ۋ���O�����x�y����)��"��g���n�ĸ�~������#rD�S�wGD.� ��-�� �$�OD8��$��F��]���#�(�E��|��
PN%?��@Exc{�?$�%9K<[�a���u n���6)�b�H{���B� ߀@��K��#�J�+�ށ�*�{#RXZ�����<A���r~¡�wĳ��}
��I>^oG(=\%�G�e�}�R=��.l���X�8m㵚�Y���G�=FCP����&,��� w�rL��u�"�[Iŏn�n7�빔��vv�`������|B��Jj��m&�5)�ga�fĻ+��� �c}]~I��a�߂�P(�ײ�|K��{Ɏ�;7�*J��2������CP��5��=�ZR���'�="�]�rjC��/�V�u�$J��cCΘ3L+'~� Mq�k]D،P������1��7D�4�@e�x�{`u`��anuߡ�=ڏ����/�U�P���p�ZS�)�v��� d%��Zo�>�%ۧ0#m(�ۖ��X���ӣ�x��V_oK}�$ik�����-�
�&
Ux���' )��[�)���`z	���[?��Y���:�;\QJB��ơ�1�a'��O���_�b�崘��<
02.�7�,���~��]n95�3���K�}|	�3˥!0B8)��K�����_��5Ϫ���b�$?}'�����q�� �f3���M�B�An���fJ~�K&|f%D����Kv�0GE@��y�$�����R��R�8F!�f�{���Ƿ���}��������3_��W�a�'¶��\lV0��۟#K��߬ՠ��/~ԁ��m���Y��*W��ʮ��TnxO��c�q�ǰ>�в���9t���..ߔ��s���p���C[���[C�|ov�.墓�B,HJl,7A4�pE��5�a�gԹ/�]qT��˒ ƑBKk��fbR���
�����j1�eh,~�����}���mn)Y���c�(ሚԯ̲�� ��El��z��RQP:�	��>��e;B���|���?$����g<�7j4���C""�,��Z�Hp�f�|�l����^l��{S�@ym��������["��-(6� �Yv�+Wp��zo��"�ñT���U����V1-�*���ٵ����5�l�]�ZY�-!�}�ډ�^[f�E`j����Êp]&{��w�z9%Y��o����w��x�b���"+
��\������W��3��T��b�h\�H��>�%�t�ee�����{�9�ԃ0�z��0p8�;]j��d�)ё��`F&�v�~l��%E̅��Og�Pnn��4�S�(g{^�g�p�f��	7�%�-��Y�U����*���2��(Ku�n@rw�P��|�ww��i���C��`��R�'����ܧ��<��'�`���u[΋�z�ʳ��B�*�q��6^�z�{���'ŅdD)��y7�_��.S>��+��o|*�\<�q�7�P�ҽ��2�Q �\����k�d�ک�6U��Q���f��%l}��Pi���h?j(+υ��\���~�\p�W+p�=�@�C_�Q�v�|V,��rݮB�]���g��Ax��'b����d$	���7]����!HZӜ��͈��ã�U�N)Mkq�l:_1���ުb��Eh$k�~Z��C5����]o��l�X�o.��J��iK�p0�}6M�<�	��oI-%=��\`���=M~� m�����RWk��W��b��ѵ����f���ʐ+�Xz�+s"���'�fT��
K��֖3+�Y0�F���v����<��(�17�S�H�lL����jk-3�� ���\�������@&�f�r��Σ6F�~؛aNuE��@$���(�Z\�S�Gu��\a���a���g�֐��.����������X~�0l-�+:��X<`X/��E�F}�\��S�e撆MʶF+��'�x��<���kI�9In1h�
aO����0��1��ݘ�<lF��0�����39~����jb�_�$�\Q�#U5́��$*�S���I�� ���0�1]�䋨_-_��tOE�A�Dh��`�u�>�"e��P�x�~���^���-�ӱ{sb~ZIgFXiZ묕�����2�X�s)�A-TB�P�3����rCʐUS=}2%�`i��ƑP���Y�k��%���Q�`�DH�Xu�[�)L���Dg���X�"O�o$�rQ�T��}�/���;��|r$�ُgI�5[�����'�>�os��b�%^V�.�WSTd��Զ��#:�nOe��Ր�ID�g���dZ;mD"�t���&P�_�.Gu�i*���ju���;ؔ����Յ�5Mͯ�pT۝;F*7���f߶�|��~���<Ju�֚�p"�>�<���F��{D�q���א)S0�+�/�xc�Y9��ezisJ汞/ەV6�i$�s�X�������p�����^����ؼ���N�-��@\��3?5�����C˻�1��u��l�8� �Y�R{ar6'���]�d���u(���ʆPr25��X��B���R�O6�R��h݃�Vz>��f�M�! ��/_�sO��-�',	&u���*�O�9���/ݎ�xf�6(�UGzv��fN�yO����g��wx\���� �zt��Z�>]R�e������q7D�S~i����~�#r��H]�Z�kc��^�J�|{�ma �ܦ��O a�ao9v��գ����� ��v�C�����8�v�Be�� �,������.�i��P\\c�\�>�;��m$z�ED�Uw
����~:�,����K���l���(l� ���d��ȁZw�w�#jxj��s%=�BZ�q,D3��̼s\�m!z:���YLv�}��^8>E�~I��]Ԟ]c@;�?!��}��ͮ@���m�ʖ���L���μ��6�h���n�A`>�X ����N�GR��;n�t5�g�ֳ֙}�O��q<ޏmlwU��@�d�:f��
C�3�$oL�I��>G�pn���j����8n��jJ��`v{k��W�����ʏ�O���	�<��,i>L��!�֝�yC�:�YQKO����Yl�Q�D	sN|=t�j�GK�9�pq�� lV���j����o9�2wkn�ྩ�n#B�Nqԍ���O��#�'|��O��K��،����w�H�������f�����dA��e^�\�q�oDRx�@��9G���>�$W_.L&�yk��}�ʫ�f�
�����%��X���_�iJ�P�\׽yQyD�h��iE4��Oܙ�s�@3���Q�!�v��C ��PոPGنA[Ҭ���������$~<'x	ҥ��z&�2�><͵�oO�B�!Lw쑢{X��vSzrwA��\U5�R�-��L|H����(��!�=s�k偦Z�V�Dո���'��Ĕ9A�%��0D(�6����p?w2������y�|.y�꫰5\�� "��ȕ�S�l���{Z�~#*0!�!��N��q����L�J�D��sHAH�d� a�U�Y�q��R��t`Y�
[����"�,Z��:��34��2���������9r2�k�k)A=�)������Ӟ�+��K��%Af]�u+�V�ܟ`y�8a(x����2�Uw�ϟ�m?�׸�#�)���Z8�Yf	��h�|[����2�\�nX2�Nٺ�p}2��e�ɀ'c��s)l�/U�X���� �l���O�)��U�6��$��A���M��[��t�>z��a�j$^�Ȟ�e�L��oz�E\-�JԀ��r9��Co��-��':ܺ��e��>�h��p��60s��O�>��!�btG
own�� ����r�:��A(ê�7ƀc����מ������#:�w�Kt��lN�[�xiNY�9|����o"��'2�,��E\���v5 ���'"�߁i�3D���(NLf�b,��B�h���/�� �'z���Tw%�<}�й�h81O#ĵK��$�J�J�k��-�� ^Y���]W��[\���v�<n�0?MP`��c2�T�� �QI�UQ�\B�N��d��E[�����z���2<��@�t	�N���:?\�sʎ�oI\,��ӛ�6���e*$(���v�� Ʉn���kBʇB�Q/?˪�llV��1�!3�v|�W,l
~��s�u��.�-�>�m��V��Z��<X��������)�o�W�>jq~�Za`o!0Δ	�W��FR�����|�V���$5[�J݃�g/	�Dnmt��uN�HR!ؒ�n���3��:_��Л������^f�����A5B���L	Q��ȧ���/K�P�I����Z�;_�J� ����{wh�;�^
���{�ƘhcA�4|= �[.�w���}1.x�o��L��xt�qO?����!���z8�I�I���t*�A�h����R��0b��۱ԡ�6ϜZ2���'�C� p.iM<�\zVU����^�)}(�X�M9^���W��QI�73҅N?<�5o�3u���1�Ѝ�ﰖ��.W�Y���g
�p����\+���%�C��wvQ`���Ś�
g$�r��S]�����ǺW�KԷ��號p���˕O���k�^˴�Kέ�2Ά�C��Bx�[T��8<��	�C��"��i�7>�AG�,��t�:}��N1e-,�iV����%�^y�$Ǆ>����N24��V2���i3�x�t�B��1�>~�����3jXc�!Ց:�4�����K�GǟQ����չ0P�q�ŤVc;����X�[m[����آ��Ւm �����.ݝdeS5ɠ�k5��O��V�^JM�rI�l��ʑ1j�]��@H#]U��z���l;�%����q����,�/�����u�dPSC)4/��l� A��u����-(/T�$+�*G�烫?�s<��_,#߭Ci>��Ǳ%GZww�Cы���������ca`.�wko����;�[�����r9���.b
�j�D⋓��Q�c��l����.����<w�^0$��������
�egrKUm�\9��Oz
t䟺Ru�0AT����^�?|��6Izs+�ÄS�!%���}C�] dq{�ڋ�i����՘�7(�!�r\tꙭ�KcI޾c�T��Z�
�T��Î�f-���̈u�Ҫ��S�!��W�#d��b�L�{/�i-=�$������"�W!Y�&�vQ�x�!Յ�`kt��z�i� E;���nJ��iN�'i#�)�8����^Oy��D�y ���Mzf݄f��]�4r�CPc�
��L�p����9Ӓ3�r�CDy13��������S�w��<T�#�D�m�*���r�a]�D"y7P��L�JI	6Z&�.��!��~L���%p}w����E#o؋�Ú��^G�'��L��t-�V��"�L6���TZ��c��Lǲ��g�o���U�E���7�oZ��ۉ+$N��Ĵ�%e��$0y-m/Jg�S�2(@t"U����@�(�"��,���	��?~��a�հ����/�I^����bdL#��)!X�{.턡�:��z}�����\㳋a���M3�;!*2�i;g���G#6�/������=�ի���#I>g+�C���|⺳���R� -X��0�n܏si����#;��Nܯf��^�x�ǖ/aP��2���$K�`��8��*Z����4f| ��*�y���rtsb�tU��'���t�c�c"�������_�4V�"/t��k�\"L/���i�A���u�x�M=�402�w�D�cQ��d�D��}ˊX�"�v��l㐓��J Y<��� z����`��db���o�O�� ��f�	�Rk��w���̄�H�/)�6*v�Tj�$��R�H�.V��Z���=����xu񳺳��,��$�ܘ%��N��`�e7'P/v�����I��ӣ Qɱ#.����&/�����\Y�bX�H�T�}�V��V<-.=�Tx���Y�.�#? b�S��,�%�[D!k�{�l���W�֌y�
7��	b�X�ݽ��h��͢���sI����uL���*�^��م^�dc��jo�9����O��Q�A��{�x��ٻ`:1��\��e�A;?�k�F]4y��q��{��x����wR��-������C���L���Ѫ�v;�Ǡ��N7RS�H�,����#���Y{��{!(��ߺ_�4�p-S���R��P�c��I���x/fdv��ˑ"�R��o���8aګG��q�P�I'�'�G%�ט��Gl'A&��*�ټ2�J�6����PvV���d��N�!�LꉵN�������߸����U�_�ǶdbM��a��'!�2�E�J�1���O�S�F�N��d*J~��o@aJ���?���mB8s>B9�R2u�5�_�'����5��3kzD�/4��/al�A;Z�/�h��C�1���f�oYz�o�zC�K�O�l�� �l� ���ҕ�C�>�/;�W[6l��c��� U��dgu���w��f��5#��ϝae�4��]������`�#�Y�P$��{�?�����iQ�=y�]�����=M��A���͠6�&`�=���m�}�K��a!�mZ�
����Fh\?�3.���};d8��u�m��EQ��sL'�J�O�9L]�m��!?�^:�L�U8~bi��Wq&�{����]̵.�2���M6L���)}.�����U?Z�,r6�����B#�D�Ϟ�@�� �,��l!�!���&/��{�wȳ�`셉�W����+t-T%d4A�wB�����M���z�5�GwT[���.�z|-Η*��nJ*����7�""gE�XV,$�2���0(�H�t�[�~_��6@%��LX0yh���� ��RR?^�z����1C�늸��L��T^2{-�p���߿gq���!��hǖ|n�c7�����q;���kS�����k�І� ���WX~�ջT�;k�e�����c���=T!5���f�G���%�-T0��9	�X���Fa�v?~��II^�b�㜨qaA�+�n/X���Lv	�Ϳ)pXtR,C�� ���hNЫ��7�A�G�=�yI�ɢT#z��x��X�P�$$5�ٙ���&tҏx��͉C�[�H ����6:i��i�-�!6R��R�A@sEQ�ɡ���*��V"
��&/��('WQH�� "�6:]�R�Fi�m� �.��d{rо�P͛�ua��a���e����P ��?��B2���lsW���g���gxZ߶���Ę��Bt���ݥKj;�q1EgC��#�/�d��˧��;�'��������2�
��Nx��_ѓΦ�����.��k��J�Uzz��Q�)���s�,� �ht_L:vp���6�ò5��uE����������y���;L�m` ۙ�>���u=��_��c�T8-s���X~�Y���4�V��R��p�{�lci��:�B�NCT_G�c�:����[u���
H��[�Y�P�����*$Qt��Y&�K��
��b�����Z$J�/#b�N7ѱ^.;��x4h�(�e�Q n��S5n��r�y�i�9��I���%S�>�5�(]������rۂ�m���3I+ʱ^�w1�
z��;���W8���i7;/�&�W9�<�99S�����%Z*���hr붪�><Z�m�;.�Ă}٣�`=o��vth�h#.(֢���O*�FAN��m(�S�!��I�Jr��h�1
k�������ی��-����
0�!�OG��`D�3J��V�����巨ݝU~�b���A~F�&��AO̢ �K�,Q�%���<Y㋠�+5��r�!4k|(I���ֵu�,^�f4�~*תּen�p�<5�;Z��p����)u���b���Pf��i<SR�`ŝu���+x%t+b6_����X�oy{���+�d����q�H��5p�ِE&O]W$����nۡ��7�s����5S�Y�iy�s�|>�ވ��J��>}����8#��r��r��^@�^3)���rԂAǿ�M0×�	z��*��,t
ÅA][s�W�J�9�n�&*�H�SX�ɖ�^��v�H��t�JM�[�:aW�V-��Ek{�,�4�)
���[p�L$P�U����\͢�D����9y�؎�CrD�
��)3�����6��~��ܘ�A=��9WUʧ�?���VGy1Y�[K�n���X��
fzG��>�,��F����K~��"&U�Po�TQn5����U�0���Z1�D4�=+f͋.>��ip�{����D��8�쥞��]���pX�d�V��f;��̍w)�n��f���5�L����� R�~��
��zn�S��>���Lji��4b`\5Y�zàǦ�8[���'C%�U8;5�r���< ����R49��P��1�_Q�sY��b���l�ISv=�m
eR����A�������I�ҫ���eRa�� 7�Hչ�;N��7ٔ{������H�}��"�jǖˏ�x���_)`��p����.H,�y8�/��u"~yn�6�h03q�e��}�3�Vv�����m�X �N�L��vFӗ�/���n4�n������R��ږ�+���ܑ��s�,�l�-��6��3���;lj��Z~	����=��p����O��*�,nV�g���
G��\rP��?����Ϲ[�;�P�&�Oy�a���^�B��K*)p��r}���Ŋ#"�
�L��o�G���<��23Z�-r�o�� Y�J��11�%�S��:��yYmH��!���<h��+Bm��L��P�"�L@��^9��/���_�ц	����,�TY��,M==ĸrs�5U�B�Fѽ`S�
X9��kfӺL�goHˠ����x��<�(�gw� �6��jw�t����z�G���6�I$91!���ł��iPr9�� �?��U8< )��&|@S��f犺�C/��w�)��=�Fn�j$N�Z9�vK��8�n!0�s�>�QB����̯�8��ez1��3p�l���?g�i�'-���n\^��Ӽ���ءߠ���g�[@�����X>�2��s:��>7m�YM�~����v��ؼw���5��[��40:6�理؟=Mӹ�W�Um��qxu�dW�Oߓkݍ�C��k� ~��1mT�w䑬����y�8cˬH�vKf_��8��
�z���*Kf<kHMo�ldL�1�t�_����;>`x+�+�3ɯ�B�n��?;Y����D��#T纒Y˗��xH_d�Z�%βጰ����F�K��;���G��;��,��*�7���ՙ�n'�4�Ifk�Ǧ��p~�I�[-@�z ��ƻ�7�����������YN���܅eC� �Z5����\�sMڡ_��͢E-՞���s|g�x�O�����ŤT�5l{���N��f�h�u��?�㴢�7���fڡ�<����aZ.ζ�k�7J���*�'"�u�~��>3IUym}Le�c�9���6KYh#V��g@>�~[^��^ʦ�y���%�"�H��ֵ`�F�W�V$I���8,�Ŵ`�s�eR\�*�Ҋ�"^�2 ʰx�SӟZ_,�����ULO�]��>h�@��V����w����}��7�%�.y.��m�?z��7z��w������bN�����IE �d�2�xH�[������H\d�m]7���}E]������s.AN�����rd�GG�	 5M9�'�4X���{�(A߼����X��n,����ԯ�l�/�8;��-L^_��È�1��?�����Tkv�Zs��<=r�J+x�߹>km�ʸ~NZ"јSw�n��٣Q��"+��rDzB�� x�V��ӗ �֓�V[���X[�A3�WEb9�6Kރ��'���o����� 	�ɞw�l�<�
]����|7�m��
�[+���r.��fsΆ(b�=�<�13ƺjc��T՚���e��"�� ��V��8J����T����m:��� �ʸ��]���	
��'=��l���ɇ%9b�^��U5�1�(\W�x@x4o��������:���l�:��"5
������Wmu�.2�D/�5�ų0N�cNR�=T)6�֬$Ԛ�ݲ+8���X�98jQ"	����}�.P#'R�0�\!��w9�!;��xME��(K�%6.Y�g��=4"ӰtQau��dU �A4,��GF�5��^w`?��7�����gӟu徿�tW}���i�(�QD�������2����pq�Y�m�E��[�
׬4���فNh��.�Ŧ��6u�旊��tr���aQ/�W���'+�Q��ܮ�Q>)[��G���ď_���&C�z�	�)w�g0��/��>)*j����G��
~�b��꩹!��q��f�xd���d� ,G����a�@L��:�F�ild.
%@���)H�Q�rEt<�����1��('+L����Oө�QG1?�^��@e���_U�ܝ4ӗ��Tړ�v �
%���P�&T6�w*d��Q��8��o��z�U��n'ߢ2/��\�kU�,֏����)d��ħx&K%P�"�6ġf��Ю�ײt�d�����';L�S������1����(���L夜5������x�-nmz|F��P�H��=�Wz%�8��L���-ءsݰUG�O�����H%uzk����j�F(�ep&a��s*^
?�E��}M#�uaxE�rV������
O{{�9)'����$؂��]9�����k�(����>�N�btR5Q.Qi�C �]��Co%�DKkU'�:Ual]_ӹ�A��U�K��lz�I#-Q%�0��o��������$��U�� ������$�1H�QY�Zv,�3�x���9�Ժ��B@��,M=�&�?&tZ��Z�m�G���.�&�c���x�����FJ#�߶ [\��"6����tZ�ҭ�|ݩ'X��6zz�+}�|U��W�?Bݜ����/�X��z]'������Q#�_�A�~� VF!�:�$�ImF��;��K'<��6UuR��)Ϗ�К&;v�._>�l��]��lIH7��MR�����7�����M2��Ö�����=o:.ɮWI������{yA���L�}�%f�ΕY�l~m~,~��o͈^��-����sl���Q��!��`�+ż�Uy��!����t�ڀӧVj��h_z�yWW�{��)�-7�i��g�����E9}��:e0���;kM~�{��l[�G����Ӣ"�8�."$l�|����L�,����^��?NʳR��w�o�.�S�q�Ly�]�_��k\�Ŵ=]�+�F������xW#�3��EX}��hE<Q6F�,�s`�U��s_Dp봸��g���D��3
� �/��j ��s����A�A�0,�OZ�u�k�k��ڽ�����ʜ�u�>�v�)>Z�ъ���WU�7�^y/��fq�a�VB��ʺg�����}�`L����o$�Z�{���Wq�+���UMm&z��Hq��ǴՔ��cx�@/�K!(8j��  �/pJQ��͝�Z\�����d��h4���._�������;9��=�r�K�>�D��ek<2�y8�'��fo�>�8�vRӡ�����N� 4�cr\�S�3E
��G���C���* e{	�ҟ˵�5�uDfG�S}{R l�׫��We�����M�oe�4
�+��N���$>_:>[�) ������|B��*��ْ5Eb��`!��eY����;ܟ�Y�b��h,#�f'8y��1��\�,Trd��q�+�@��
#�_�pmv!�w3H�R���+o��c=E����l�������:��`�����6n~E0�	Q��nS��/��r"Ƶ8��x����6*�Ɖ�,n;B�VwY�ô�>�_~��P��?�˸���=�����t����3�8���H��s�\d!�u���*C�De§Y{mm�5���Z Ct��xp%V�x�]7~� 	�=��Bq�*��H�KlD���;�;M���W)��d?N�-��v����X�R`|&OV'=/�	��¦��`����;>P�r�5���DW�����1��e���iT�s<��aT������~��m�9J�����8�u@
*c��/x���-�H��ǟ�GK1��1��Ҷ��;7w-AQ�Hs4,*l=8��̛���⒳�,��4�̼U�J��i��cfs��B�_�[��Ԛ���ê��VE
�-{�oew��`F�z�1^EK\�_@����6���:�7ڪ^^����D*�j2+�<n/1�ܘ�e��������FJ�\�7�yE�5�M����X�0�03Ӻ�Lӛ�d�O�ď&���w�h,�,���p��J��M���7Igj�tم�י�(���Lg\~��x�wfoiፋ��)�!k
z�q�����"Z��
#<��kI.��S�K	#����e#&v9�qq�4vZqhx�uUϧ* \)�,k+��Va�ߨ�`i�g�NŚ�+��i�������¥ � �H��c��"��5�>�[�o�������e�s���P�斬��V��q��	�22:�����Z��i���Z�%۶+�q����,����˳N��3!WYD; ���_B�@���ذy���8��q0PB�]�sm"[��{���od������A@�IC�����#y��1H�o���M���"_�Bӂk�)`yZח#��	��U���fN7.����$9ܳ�E=�{?����Mk�Oo8��䭠�㹩ե��u@jZ*�E��5��Yq�����V12ܾ2p�CV�Q���U���$JǑ���Z 	]��"�K��{2{�E�9����������%Y@F"���❦�1�c�~��v�bD���;�.�m2h Om;V��-�ْ�=ؘ�W&������ {ח#��^\�T��m}&m��7f��sa��u�J�r!��h�.���c�)�U<"MAy%F���*�Z���1�@������o�[;D�����o/!(y�uy��+4f�~�Lck+,H�|7zⰩ�>��դ9��4����YIz$1�R]���A�kk�}y��xp��?�,5`(p�x��6)N�u�W^����Ԅ�`�`Er�=�bEl������p��e�?�!0,�_�x���ʸ��٢�Y�q�|L�*���o��Ju���^A
u%��>�{N��׭��=t���4��mO?M�չ��P�4{�e�S%/W�ɛMg�nK��d�)�Ъ��f8��|O7���ym�	M����A�4����^8�&^66�*�'��c�9�7��d�+7�[��H���KV)�Z6��+3�KbΎ���ZҾ`��[0虪��D}��Y�&&+�e��A��\!,\�~�v~��rX`�Ju�')���cAx.���Ov^�xo�>��B���H��KP3"�fSb	^��b��!�2چ)Zy�4�:?�ݽ�1?yT ���ҪȝJ�Ӊx?n-U��0i!8�6��#F��y�(�	����ڥa��j@��d��P}~m��E��E&elH޻��f:pq��?|�闄_�
��[;�T�^Xa)��Ud�9�,p|��蠡}�l�_�Ҟ��O��8���o�~��67�Iڱݣ������Q_�����O���>1P/�kA5;ʡWF� $�C�O�`��>���h�tl�XB�d#��4��C��;�!��� gMVB�_<����j�Ԗ���T�����kRs����x=R4Zpa���=;Uq�[����7�u� ;
����4�G|燒��%���f>M>��gN��*<��d&��S +�e���x(�xJ��oUIa6�����Ҙ�5�)#�9�b)�=�K��	x!�R��F�SPF��[��,&��V���7�[
v4A��t��ic��3�J){a`�gsjQῼ;��e��SF��
`e-c���ģh	�
H��]A"ϧ�x��m��ca���B��3P�\�jE�@ǟ�5z����cÈ>�V������{���U%����vO��C�~�>�U�1b��O�=vD�:�6c�ϼ0�����7@�����cy�*�g��6 T���7�)4�����V�,8�e� ���g���l�l=��e�G�}
��{���2�4���+����1j���0>g���%���
�] $�YD���|g���*�՜^��Q%$���t�.\��鳳��8��C����SUjF?��������h#t��	�ri��%%�_9ޟ�G�	[� �����Yؗ�,��KW���K���;�� ��^W�������A� 86jQ@W��@w��;Ԕ��[+*;��F��V�?w R*��P��}�)N��1)Hj�C�u?�D:g��"o�g
M����r�6Y��WC4���47���ϕNpy����hd�-m�=U�~r�~��+`�YF���Cq�]qr��+�r����'�'��#��7Hj� O_�,�{�@��}��`p#E���3�4���I*H!z����ǌ�:�MMV�G�K�:{�ָ`��Y7/2޲!�dzD��MH���fu(�)�;�DZ~�v.]^�AG>�"H�חZ��ZO���Q��#��`KJ���8�z�5��ɗ�^g|��KDU��żL>+ʩ7�&�p�%��b��gVE~����[SEtP�$-���^�C'�7�����` ��ۇ��"dR?*�Eu�{"w ɾu��L2|,*E�
>���V
�i�	
�8�yaS"w��X�a�����6`�\"��E����Z�?�H�dwq�ǻ�p�^=�\Oôw�k$�f���9������_�,�?6R����I�[�kd�	�a��+���(�ij ��i�H۱�esi��D��0�=�$�v܀�1p�:�A��9p�"�]E���=�%Ȕ�0lvi�f��_g�J�a��N�{,�m?t��񗊹+k���F�y��X}�ϯ-����>��g�6�BGD m�SB���x��u�>8_HH�x��?�K�`��X�� ����B�KbTi��J&���J'b�nӡ��>�ᴍ�	C�kΈ�'bP& 5��_-0W1�wb��G�i���9�����=f�?S=n�m���l�w���Q�~����~P�\1lq17p��b�K����v�nb� ^��be\��D��ދa��y���i5}��l#(7)�3��d�R�)�#y��3�E9�3���/d1���0��7Y�F���Z����΄X�a��N����ǻ��p�?�uZ��@R��*�q�B0��b��Tb�4�6���|3��3X���G��d�h�A`�!N�W�N��$��Zv^& 4G.x��p2?��|k�Vأ)��:T��`X�xp������a]ꒃ=Z\{��~:j����{(C ;��|��:+NZ�c��&�[/%��\�@��A��֙X� (�6jVI ԝ0N6�֦�+���<G59����b}����=5W�@(��,rz�H���	)$n�Z�tƩ��18���7���s1�t�E����3LzH	����/7;��Ȋ\��̏kA�F�=����N��W.�7�[�=�l�L=vXh��AT���DL���<��SRN�)Oz��8*a�O\Zn/a}�����p_�j)����/����XO�n|���r�1��fF_pU\�\g��Y��62�A�;�F���F���\�ˉz�8�k��p%:q�r�W���M��<���Ր���.P5d������1Hx�U�1X�0;��Ë�3F��B��)o᭕
\��y�d�5wk���N�<W�Q� ���9��u��M��ae�G)�$�Q�7�R��9�E 7�8.8rFk��cP��`3ԟ�5�"|&� �BJO�f��ľݑzZ�N`]7�ރ���|�1����~�>ZR�v4�(պ��J�Cx�Rz,ߍ�G��1�J-}�J1���v8�+n��j�Ѻ}�r�ƚ�4p�4���E�����/>mui�坰��a/�&[?�z=��Cí�vjL�ޠs��7z�[�[��U7�s����y ��Ҁn���!k­19kOᣨZ��BUq�}/Mk���]s�hX���P��v�5�,Bn~�[G5�x�h��6�~U!��41N CFU���A♓�T����uUTg0;�+�L2��[}w�".�ӂ�t]��۞N^�^Y	�oND�@��Z��dԿ�9d@@�UqkJ8ȳ9ˬDx����%�:�UiA̧�$��sj�޹;�B&�QLS4*e6|�QD�����ӂPٚd�_�0��.�"iRy���^g?��FB��R���=��Gu�<�{���cG�oa����{;�������FI2��X�a��iW����dJ���]-��h8�i�O�܅�[r�6ʶ0���x��ӆ!{b>K�GG��z�~��]b�Izy���l��7�85�����g)��E�UM)�a�5i)Dt}:��;%+~]�+,����+�R Pz&�Ssr��g��GU=���zn�C���Mw2�`5��@C"YL���``���+�o����A������I?�b9ɼ;�^6��!/|�Qj�G��Y�P:AE��@^��Vq�#9��+8{�Q�8�ɮ;X�+@�� �l���7ne�g5!)�y�R�t!��4f��Ծڮ!��g���f��zM��zvϖ�U�����WB`�Wf1v���浲�4D����Z2�;WB�����l�ji��K��k����T���Kt�VaS{��b��W����ja�3{�`3%և�R��)��`����B��Nr�;]~�����OY�KG������{R%0���*�t��G�(�֬@ܓ� �_��	ro\�d��P�m��@�+�K@�4�������A&]�!fzMGo FǓ�OdS���`��� �|;��N͛
�lʠl��z=|�̓�Kh.�6��a�/�����~l��h�X��*�-U�S^=��2rs)MB��⁝X��*�K��ql�Nꦩ@TEs�v'9�F	-�@ڠ�g>��ў�9"O#�����O�.�3G4�6�h�tG�����i���/�M�#C	`X���=�����n�%��e��5m�{�|ش�5	�N��omi��K��9��
� ~��!����x����bS=Ʀ�3"d-vC�{"�\�?a���˵���~9����{u��N(�U"����^��U+����yP�Ԣp��,��n��eW�J�?�W�8!0�E�]�0tt���e�-k��E�?�⤘}�C�!����ƙ�8��+^$��zGF����l��cf v�����c�ئ�"�Y�$}#������� {�R�$��5���P�E��(Vm�~�����9��@�%<���}��L�t �<�6��[����O�-.�ɴ`�s߀�Ұ����ʁ�.�;<��LQn���@��� @e�Q�E��@{��{}I���j��N�d	���q-�_�jM�����zy6m�w��	[ҧ�d۔�3='tjRN�?wA���rQ����0�c%km�.��@O:շ�Cz�d��{��9v����_kr��`�{^7� ��#��А��M����d��u�'30��mۗ�����BI�������-*�w�w���V�?����h~2o��#�yA���Mb����$2q ��y|��M�u�A��#T�1�{oDk���&��B�&3ѝC�-�c��*�����P�R�9$죄����h�}}�_x���n��\��ip9L��ц̦��Os =�dh��P�+��u'�?eB�6_��\|��yŝ���z&��o�7��wM��j<A���9O%�#Ϻ��:�����^�>,nl��d�� �H�.`� P�p�4X$��(�P�]0���� n��M�d��-+P�o��b��K�4	�'���L�F[¬9*d@�bo�����&|���;*�'lH5(��<f��E�g/׆�βiU�ed���[ J5R����q�bۉ�m��H�r���	�'��γ�1?�!��i�b����:��J�^����HgROwC4&_W]�7��Z�Ov-Q'�;�O�0��hո�*��Z�?�{7H�mq6H|�ĭ�)�7؎�P��@"q�W��E�I�Ǿ�$�`��:t��@�lml��\%_eI񯙢c�'&_��(�ڕr��y�`?i�ዃye	��4�-��;�uޡ����`\��nD��A7�4v� 1FKQK��4������Y����M2����y�'�U�L�tj�*��w�ړj��3�ѻb<2�K��s��	Z�+f�������V�&MZ��,̚N�����_�EE�^�ps��4W�#1O4wl�ӭ	5�S����I�\����9��Fd��U
3�Qהv������P/*�������h��Zn��P��P"%��w�ݪ����@P��5*�$J��Y���C7%bO���c���.#�G�"�(a��8�?�5�ԅ=\�p^���Df�P��}�H�נ$�r=�=����L�a�f�����Kt��&͝�q�{|&����-����%��DM:�h����Y0	
s��|�n��+.#�_�g�P5���l{7P��e�����_�!C`HĞ�?����ĕ�L6zo2�d�w�R8� �b����
R�˚Y��a5BQЈ�z⋚s�
�l~1�����zx�ڥp#�P�1pw_��d��+ϋ�|�z���SlF�kOk���Pw�����ksؽ�iFf�Y���Fo�I�W��'�Q`��ܾz���6��ƺq5P�X�`����nk��L�)(�Ì;\ק�N�ێJENJ4���q�{/��=���$R�H�j������K�n��l�'�+q�:�����7w1V���cv\�]{����%4��
�	�F��*S���[��сV�v
�N��f�G�y�f���	���6�(�z�6��Jt#&-�5��S��߇�ԥǽ�l���: =��п�/	.BM�q�֒n�U���g�����G�c��'�.��Ne����Q���1�i�����p�^��Eam�T7Arզ���`W�9u�l��-y�ψ�?�l,(1wZt����}������d����-Xc�����k����:x��v��s�������ܶ)�(�H#1�K�9J�-�.�wΗ����D�{�N�k�G����׃�����[�Y"2�.����G��F�sݽ�R��ݮ=���q� ��;�r���jXe!
�[����[.7'���⒜̩p(�\�'����Eb�������eZ�w	A�EfT8��/C����]�E~���Grx3�4�����L2\�H����nqct��'�����z#�_Hj�)�_G�Y�����ɵ�-_h�P1����.d5�����~���EH[���L�pn��J�jXm�@,�y2.�W}�!���RS������b�nթм�ޕG��ј�q�LZTOg2����M����ܞE�g�!�[�����8[dV(����Z�_f.
&i���R����¾�xG\p9�Q�AU�1N���+�G��}Μ�`�0��~/rb��9ZU��]nL�{�?g`������t��O��vp�J�>b�y���*��f�lo�3P+7��^y/���Υ\Jd.R��w������K��.R���=b����.�-����ɚP���u�yM3i�H��hO�@�p"���֫&͆�b�J4���6���x�k
*N׆��b�)����N��è���k4u��(2j�H�r��*��0��[r��!$��W1�����յ���]��F��I��R�o�+o]��O£d�#;!6�aL�%�(�"�������/n����=�z���gP�H1J����Z�[�A��w-�Mɾ^4)��+W�����O��`����;���Nx\d�L�AX>`�����艥@LYj!(��3���{o�S�44�!"�;�]��&zBU������A�>�gM�4� v-����*���=߅�'�P��x��������h�ٲn{��SO�軖
@ʆį�$��G�Y��b�;D����Z�%�pZ�`T�ռE�,����	2�+(+�fJ�����x�3��7CSњa03-��cZ���\�;i��)՝o�П�l�׼���d�L/<�=��4i��NI,�=�.�U~BU;WYiUA�Q��-�4��h+y�����X�\
	�y[r������*�}a�2��³Ř�GR3� 8q}~m[��̆�9/(9tm�(IȾ|����s�	T.V��j����e��B�d�)Γ	!�ܯ��D�ZH^�zu��{� 0�[����L�Δ -�V�L�.�>HW0;�K���n����P%�z���.;9b��k�rQ�d�ĳ�͋����ϴ��nG]�u���̯(ڲ��5`� �$c�L��g��x$�j�d�n�0���������D�6�˨�9�����f���#��;�
ZְNSr���7^#��u�Q*Qtp/��9#~c�y@�*�d��`�)�%����.M���|a�M+���.�ٕ"+4�h�����m�U/��nۙXcD�4��6������/ܾ�5NJ�뵘?#A��c�4EO��A�ItVSY���-f_�[*�I�d.�6�Y������q�sb^n���~�Y<�~��$��Y���a�:���Y�\�9��C�ӛ�@��.)�q������Vhr&6\\E��
0i��Ĳ?�Ϗδ��7�$���)�Ê!�\�&�����*q����bezb�
�h��n��X�/;�4���x��;V~�2״���F�"'a�7��U�����N--M&`�l�H�
�:h.[�-��/�poAC��TMשiR�8�����e:bp\�%9����N�8�p�`/��Җ<�-�/�� ���'���>��ߢ�(3�N�o!ڑ{�H�C�}
�+?
�"���v�r� ��}-\Pl=�2fM�X�!��b��WM� �ay�y_j�/L��p���9����fdl��2K�}(x�=/7Z���/�$�r���_�k�������*W�+t��i�{ˑÔoV�o���;�t���.��H���D����Ȣ�_����LN�cF/{[��䰐�� �c�]��qү�?T��x��S����5���n4��b�k���Z�Z�q!�eˆ��mG8 �I�'�\s�T6]�<̐K��eH���짉��s}���>�8`P�^�,*���-�-��4"��R'A��du~,��vC�Y?~�8G�@�8{+F�"���Z� w���	ӛ<ܚ#6Dh8d�C��<��O�mh^��Hq�'n��՘�O�FHdS�ʝw���6��O��T�X[Ƕ+�-Y;��Q4*���jW*?�-�����H����di��R�A�������;�86����H�7��aA��P�����L�||-�95��ھ���F)���ʴ5��E�X��,�SH���U�.��wƘ���N���D\[b��Y�Y�`zlYJVf��K+���+�hW��A����jJ߾����jPFp����+���Y1A��7��:'�n���YB�$敶g�=`L?
����ƀ�2rv4&�$�O���(��/�����س�J���@���+�����w�G�Y�g�i�W��z�ڑ5;���r�X�e@�퐷4Y�"�\�`S�32h���Zr����L!��i�~�~F�f�0:׎�4\`3�W,����-����� 8w�e�c,<scc���w~P�7��<���
�������He��Ҫ_vz���<7w��~�&(b�h��9������6k��<2��:�erg�[����SW�U��a��A�YÑ����?mڐ�N��#H��gƛ��~�IX%�<�<���j9M�S�g �����$���"W�(�Dd�2d����ݨ���A�ȝ�v-�TG_�(͹L2��4��P�������H\i`
cj�\���P�����P�ho����7�pG����%�1�ْc�v��#�׮� o������qjF�\<��^�/��smbLS��L ��{����/>��.#S�� ��ڱ�;wFKMR���ԣ����0�N~�����x���H:���3a�Ϲ��&�F@YWr��#��SY��Gv�J?g:������Z��DC��d�;_��n�������x�l�
�ղ�m�Ħc/���������k�۹�}���C�Hi`����Z���3>� j:g�N[�%�".r����s�!ڳ�N�W��*���5�ҭpڟmi
we#���^L�eÉO��#d����֣��|h7�o��"���U���{Q[�g*嗕��$g#�e�d_JLM�88��Yٌ�#�i��j���������� �(��i�~+X�� ��&�:-��� ŋ4�B��2";M�yu�V8��tE%CDC w����E�g�eڋ��VUÎ/|��.ߝ�!�C,Hl�����f�Nh>��gr�;^;M$��,sf9�u2�8��J��8Y�)@�F�.b�|��0���\G"�܋�%�C�e&ZY�̉���h���}/�f����`YXU�@`s���`͠�OM����K���#��Z�48	�dm���
dt豟hj�>K})5���ٍ�T�'�)I�2��jjKq��`}W�n�O4t�*6������f'����������3�uܛ�(���ࣔ�����L�*<�	@u �:����z��OA{�CT �9:��P�	��}�8^ߥ�I1�z�r��y��Syn�^{|��G��)~�LM�P.�K�F:�"��x���<��f:�Ll�����͑k��������
��1<ڰ	�E�E��s���[4���bX��
{��y����R6��f�X�!�6���"2����H�n��[ �oo)�Ͽ#��D���������Ȑ��S4j[B���2ؗ���J)Ax�5H	��?*��m3kp�N��L�S��kuY��'6��n�6�� ����kDQ�(�����&�ykqט�Ŵ�g�34��ȵ�%�vtwK�P���gп���l��6��Og���ݚ�&�16
����<B蠛� 魛�k�4�*�$7*�Gҍ��3܀��&q5u`�O��_8���At��}���c��`j~	Pş��kR�g�W(�IN	���_��WXG�Z��	k��o���,w��q��������+-d���t����C�X�籆��Up��Qm|�W5�i��5 ��=p�6`D���5'6����4TM�瓊�x��O�W��F>��E�g�ۮ�Ϯ�b�$���wY5�մ�g��T+>�^��1��䕷Hb�>��(��5����&��o"7.��P��(l>޻o�PY�n��-��-��6 ���<��/W��iڬ�N0�G��MQq��t�5��t�>o)�F,��:� w�ܸʓl�#ZG�l�<̪W%���"]ӧ��O�JRg2>h*4H�'X�)P:N>�ک���	���)�Pi�+���8-=�y�u���M������Vo@��Q�/�Of��L �;��צI%��R�4�tD�c�,�0/'w.K�R�<6��~����+�/Y��*��Ky9���`�&�aH�׍J�8F�)0�@���׭�����n��F�~�X���tN��d��@e�P�Yz�}��br��� �o{fG%P� �����t.J����Q8��
M<r;T��F�9a��`�G���9[���5j���e���G=�����Źq�kG�9�/}`��vr�u$����DY�)T)�*Ppx��ȫ?od�k]��f��?#��C�әs}l�[m�n�B��<��愳��1ߎuY<m��{���r?�aW����t�D LǮ��kH؋ h����^gV���ʠ��~��I����M��d���{R��]U<��
�g����9���;a�rm��	�'��,&غm�������_���̸��T�����<�����0�L�LB+*�'����AWK�e�	s�ܰ���<VT��CM~���c}�?,�bC~���ú�s�A�f���a������#۽�5|Φ�:�}%�Lf>�d��0���)E�$v�A��J��>��f?�ۺv�ˎ|�*�4�.f�Bq�?�v����l�1���[B����N�p����3&�څ�]G�k�AI�tA��tD��xKy���&��I;>ъJӽ/sA��}�����mY-	p�t��Z�@�I�,��KFӪ6��ðN¡�软 �qݍi�3<��y'���H��rN�2Uɍ�+�i5�X�Bf>���|Щ1;%�+��ŝLi�a��,��Y�f%~�H7V�l�Ľ��!ʺ�"�Ru�j?��zH����B���q5j���t7�6L��4 �SkL��xD�^9`Kv~��R���se5ȴ���%/K��%6�&i���~�!햒�P���j-�G���Cm��3Q?�����awRz�r>����]/徎i�R���e��e��ĭ���\��ꎀ��o-�+��12V�	�0άb��d0@6� +.��2]"?0>C$a§����+Y��͞���[�f�/8��A%�R�+�0L>^�n�w�![WLL�jT��k�o�E;h�$B{�sx�.�Q�:Z�g�R�p#(Q:�B�8M���.�)�"S��H�_?ݿm�2�ꀿ"��]ѡ.���0@�������SK_�SH��te���U�ʖ���[�o]���6�j�<As�Iۄ����`S,%.�1b|������)���t:?���,��ұ/�㉐�]6�Y��>D߿��?�7�^by�T��QU�������<����bQ2(qXC#��
ɁY�~����`ÁΡ�j1���E��RE�һ�$uy.!�u#f�[�xB�t�*q΢ەūf���}���]<�I����Q���c��?�^�Ļ\xݾ;)FB�[X��k�5G}ֳ&��	#�M��e:R�wk����'����]�"�s�@�8�4>>�5��	A��Ͽ���Ihd�HJ�̠����s�l9�S�r7a��QΉ!@2�0f�����u3 o��ʥ�X3�9�
*h��[! �=w���quߖ���5�  h�XmqQ��{��OvЧ��8������5���(&�2��K9��ĳ���$�T��������4�i>-LI��i®�����&%�����bUxQz˕d��]��
���>L84r0�q��z���6�'��|�k �u�p�'���lzԱ�+��{$L�sK��&�O�m'xj�#�)���\D9��I�w#�;�ma���D�o�[[ou��` �o��	��*�����'5�>/��6�Ӡ�p%�WA�"AW A8��$�5���"���<V#Kt���Hix�S��]}���O�a�o�R��+�C�5"�H�Niz��!�=mt��͚�[�n�؉Ņ���{��v{�Y��&G�*N���!.�2YD��5!� ����ć��ݨ툫,y�+�	"g����t���-4p�2�4�|Ởd�	��SeD� �MY�xZ򥔀u�����@G���������꛳���bJ0G׭��cO�2�����>"�<�����&s��ߋ���M�I��Ɛ��U|p�}a���R��ܝghDI��ǩ�5J�����J�:�|�0�H�D-*Nh�/�m��+��t���j 2��~jV�������	^�id�ĖU�{�H7p5y����,�O�v�E�Ӭ����(�I�ʠ�p!x2�E?x���f�o�6�9~��%_=��i���C�d��}�C^*�W$ۏRm��rُ"��[ԅ �v�^��7��`lv8�/9C�9�$2�DVB��_���=�܂����M6l��^:P8eN�BAb����A_��5�Z���m05'�ǡ#��3��l�?�똀j�b!��ٞxC�J��k���jPl:��K���ybK�7>n S�.��C�;F�7v��s������K�ﴸn���횖%L���Ft?3J�)E���_�����^,8ĳ�����*Q˫���J���P����>�L?�_�Y.��n�� 	bY��Eu��6�p�Q���y��ڄ;�6b��a�CzK���L|j�W2���{md�sd J��ī�cb$�LPC�P�G���|P�@�&p;7PV���/FS��1�΃�¡`��e�?�L���q������7qWP� �����eB��pH��;�����c���G�ᖶF��AHj3E�3��J�Wɸ1���紑̤p�3v��=[2z�� ��[��߈��!���Gw�8IG"኉����K��%,� ��n�W=<i,6�]v{!�R�\��123�9�����F�`H�x����M�*R��%T�0X��������Z����i�n�Fv�?��Dwػ��*}�OM&���}������{�d�$�m�Iꐈ�HV�Q��א��kp�q��/FD���v;��+���w�f��k]�����D՞#�����G7���7�5ﯶ$�;�!%Bլ2�G%W|�i�G6k��1O���gMNY�W�.����n��K�x��S���k�8<,-��N@?R�������Hy���Ҝ�o}�w���)
.�i�����R&�?X��i������:�3]���,�,F���X�)R˯y����zd?�l�0��)����C���/L{����̹;~RH+���H'��V;Z�H��5�$$ M����{�ME*���d��wt��\MOĚ�Ip��������񢬘�p�\v��@*T*��veO��2+�F�-�^2� d��!�jq�q�q����>��v%uX���Aa�H�}4P���Rܠ����V�U��������^�+�|u(V@����ĥ�JAA�^�6�&aCgn�bХ"0�x����g�؍'ϥ�����h�_����"m���4�l�������wS@��SbD���t�^��`S��.���]��X���[?��ʏX�L�> 洏�ɂ��UEDV �v�Y�f;<$��c��d�o��N ����%���r5��[����<H����$��sO�?G ~��.Bí@Z�m��J����*v=4�A7k�/��bO"O�n]v�a����0�X��LA�-}t�X���c�wcE��hS��=�@)D���ę�,ړ5�yZ���yD ��깑}�eKQ��"��0�d�w~��C���Ѳ�) Wƣ"1

9��B���g��U:���5���d�G�h�΍?3�m�r�O�h���8R�����Byw�Q.u5xU�b���yWz豹�gdq��-mU��َh��ԲN*�m���a�2	|�cK�_c�(>]�bV�JL�x��1Ƅ�+���?'�F�о�:�!2��k�!;o�r��F�tg��*M������v�f���ݑ-���?/Ex�]��!����z+7	ڭ�"� �*��u���o�aG�]/�'Τ��;25v�Ǝ�9�Asa�DX)VV�\�$f��������+�C'vv���Hr�����;�8_�-�[ /u�Dpo]�E4��ʒ�F�o���(��g�"�V�F��Te1�H�p�ߢ���bR��Ni�"�
 [��m� `^�3/PԽ�3��v+B�L��>K��ƫ�Kr��S��SO���>]X�f31p҅޻�9�ד�m��:�ӷ�E=���c��k�s^'h�50^b�\;m���[�r�Eٕ�sE��q+��x j��3~�oh��|�	�0�)�<C"T(��Ч�-�0 te�s�[�s���6�����K�Ѥש�G���Q�C��Ms,���'��b�Z="���0�&�H	du��X0�f��Y!dD7rJx;�sB�]��m���|_E���vX�,+ؿ$E�ر�d8�����j�B�ۺ�ĥ_ɍ�)A�"A�O��1� ��׀35�+@�ū>������<��i@*��O1�n�'��=-q�ܻ?���i�(s����
u���[eZ�E#�}����wnj2S� �0rͬha�J<t	Ǔcm �~��{�J��_FrcO��ea�O�XoUG��Z1Mu��K�qvI�y������K��F�o>5	g�۩��ckiZ1V�M��"��2�u�"�����^��/س��g�5b<c%�.�κ����jxԎ� 
QG'Smx?���]t�@�6ds�٤h-Bd��k�0��t#�^�Ho#W*(I���(�4�`�"&.݌�����
�:i�M���	���~'c�1��^{S~�v�h?L� ��#��7�%㯾��Ƚ=�e�bcؑ�֎����?w��j<��tbˇ
�_q��x<B�Q�;j.)�4qǍ&n%l� y�ZM��Ҋ�<Ӌw�i�%�R�Ҕ�f"��d]3��ю|���&I��E7��ʪ�T�J{p\� h�ݧ���g�jyb����M�x8�]"բ}� JG��q��S2���x׍�UJ:�U8�4"��1���tG��en�
7��炋���f�#:�� ���R���`&U� �,pc^�s��<*�˖NQ/�"x�U��`vy�������+���`���L�|�NExw��,��Ev\ǋ@m�=�?iזy��Xm$�njf�ŉ�2��D��>e�Y�IQ3��"�[��f��4@7���&5XP�Gy�ڷe��#��-y�V����:_���zA�L'5���F���}="0�a��d�)���荼x�-��^���g��=��,g��ƃ��g,��S��]���.�EFo^�����!%:h7ȅ�H�/31r�wu.ɿ�D������Y�IK��-��ݟ��j�=�F� ����qy���쯴.*l��J	���<���]�J���X�-�m��a���.	=o�\X�&1�"��^N��	esc]h�%���/���wo�aP
�o�ۻ���CeN�U�x�����-���nƕ���Y�2��_�R��o ⢬�%)�HZ�j�'��e:�D>e�p��b�6b|�O4U�?���	T�mw&(�X�^�D�� fW�1�(`Ŵ�Kc�o��!�9^Rt��_�ܫ�qH�SW�oeRTݶ|˨��#M��H�7GJ�e�ka���x"����։���RB�">�*����?�hC[�DB��?Рc�S5艻���:Z�������a���v��[�_����.��;a�5�zR&�!�ƾ�-J8�$0�'��:\ �1�1����L�ꦟ�B�;:.���u�U=�_�}ֻ�_!���X�q�J��5���/�e��iG��ݳ�z4>*�x�̷���o<��ۢ��1��,�1���P�M'X,�8Ŋ�-��ه�}���ρ����[�퓤?C;�|:��3���ap�$!hG٠��w5~$�X5��]G-<�@�VU=�XY���x{���Q��y�c`�xNW��! �)tt����I�{}� �N��8شh�r��~Y��=z,���/7{"|*����]�B'Y�^2�r.�^,��\��� ���_V�j��P�q��s0E�d�"�I������{*���������e=��\�6�ټ�#�8��mrӒ��
r�=� ,���M�<�k�(�'�t�D� ��]�<}S�������	Y%n*���V=~k~y�r�鶂6�c!�Ӱ������ۼ�fL
}��]fN]خ#�;���6�~{�nT�����o7.Z�O�xD�L���[�.���v��=�ik�!z�Y�WxZK�L¦�ѡ��&������h�����F���H���P���TG�ֈ�aˤ�_��h��"LS�eb���Cf�@�k�j�!��n~��e�(������VMwkz�����_�����cw�Q����M��i~tkZ��6Y�+1E�������c��˾�s��k�3eß=0߶�g=�0�I�x�ߕ���O��ث?v]�[�v��7Ҳ��S-��g��h��-��Ǭ_�ק٦+�W�K9>�I_������d��g+�γϊ#*�;3��$��y�A�3�V���Z�ζ�jϝ�O�����Ĵ�'#8�Ҙ���<5#~�(�,�����:Z/�L�s��@^].�� ��r}XPX7 �r������1Xn�f��XN��B��ԊZr��=��>���?k�M�m�1�%$���f�����)�9��E�5��ARJ��6xt��ؔ�z����q������zd ��k����@�2*뷋�0�g�pY���i������a8rQD#t'u�Ζ2��<Ñp&�S4U��-����;~�����(�h5��F�����	� `���������	-�=p��K=���)�ы.��k�6Ε�|�=�W����(��64'�����g������'�|�viQ��nd`���+Zڲv��<�O���N����#X��B��X0o��ԭ��V-n����{0K�Մ��`��[i��m{���O�Ʋ���m��� e-��U����<'�_bP#%T�1P���#P(���&n�[��˨c@�d��Κ���J�&�b��*o���;�~vh��^̳��`�ӊf��Cħ$R�Q�����5vh8ޤ�т���6��V#����	S�x�|�C�g3���]C"�69��Z~���\��ɻu��]:�W��D������@[�Ǚ�6�> �)^~f�M֋q_��y������De�=Hm.Iq0�d�0�:"�q��H& o%�P/�UV��v
Anӈ�#8GZ����xW.C�0��%�=��^c��F��o��fv��l�w��:�z�NR'�A"�De$�>hS��A�v�즜`cQ@�EUw�)���b��
���=K��-������Q櫀PN���x���=X������6h��zW�=��l���M�����Xa��|0�:^�����ж�*
"q����H#���D��97��G��ǈx�J��wx�j�q��W�O�[d�>�����6n6���^K�֙�]�8B��Y��m�����j�b6s1�:���,�Z�wٙ�1^�4�6�ڌŝb��c'�Y���ջ�a-���.�ڢQ�2R���,T>�������@�*ݻճ�Jβ*����2���2��v��z-�}v��.ys%��	ŗ@��!���uA[=�_H���{��eP��k��D�&��nuOHBec��zߌ��e	�d�áΤ=r������*m=
g��l��h������[�u1߽���D��-]1�tޏ�ن̶�ս�?����ݩuT��8�$���`i����ur���0�u�!�Ś�f�vSU��fjΕ��%��t`>=D��qz�q0^��:��H�%v�xj��Ud�y>Kѹy9�8�NĝX��6�� ����ف��?!��?ѡ�uG}�4�T��68p�d�xd��J���s)"��V[(@xS)X.��	|�,w��� �-���5�(?�ϖ�b��c�ʚ̝:�f�/մ�4y�h��n�&���о�B�L t9���8�v]���Q�]�gג��q�!����|_m���=3/�^�r�C���$|o�-x�o�Ɗ(�57��s%G{�B3��W�0�ou�M\6�761
�b��ɹ�l瀤�R�n��Ђ@��
s\[����+B�
s�5��s�Q��
���m�&~��]��]H��HW	�3<�v��=����'n(��qG&�{�@ ��.�+�f}��/O��vE��
��E9�:q+��4�Jy$��L��fg������jp��������I�=�g��<O�ܹ&e�J(�z;��%7Şd������'-�#Ӊ�A���d<S�4�R�D{����T8�*~͍I,��a2�+6y;<%q�6ts�l�i^浭y��,��Lɒ2,�(�~V�[O�L��W��q3�÷	Љ��G�㊘�,_/�s�D*�w��ٙ��-��)b΁u��_�<%#�R�|AV3���?qU, �.-��b:P���DW�WɾD�v�z ��s����6��\:q��
����4��3x|ۤk�w(����+�����iL �}�!"�p�-��i ��Ir�H�R��H�%V$�X��{-�"�_��ŀ$��/�z����\��r$(�m������K������)�zX��փx����j����<��d�e&؝��.��R��zhl}H��Zm=����������b4��Mdի�tt��'�z-���uF���L��HP�B����Y����$u�^O�)�$T�̸l�����-T�5��A�@�96��D�p�ԓ֜��Ne��HT񴄯�m5l1�q8�NH�ƒ4/s����q7�z�C6Ҩ�V����s�k\DU���U5ri��}כx��I)3����(�cm��~� 3����9�EO�O*�7�ݘ����.�c�ɽ\�4�=� �R���.`·�z�:t�w��F0�@Ǭ�1|m�����ބ���)�.����r�@�d��ͺ�jn�]�J-�!8U�e|���d�A���cm=�[gY�4�c�;�f7��Qx�^�n6��+���͡�g�r��vIn��������d~)�k٬o����~��Sb�p�!�u_A��mM�� UzFs[t��q���,�r�B4���p-d��27��JσbA,�m<d=v5��=;W��cj����ϤۍXϥ�!O�Z�����G���s�.�B��C�˛⢂�'��C�U�)�i������k�|���AbM�/qcj�3���^6�C���;l�E���O_���A��(�֫6�;�������I����_�(-߳��klʛ�{�Ӓਥ+�;o܌a��;s��S'�fI�~���,�~���ЉD�-Ay'A@�I���f�+�qs_�R�zd"I�$k3�?%�?s��E@ � ,���8;�"M�/���7��$��t�c�c6����/0G
VPfO
O4��R�h55��eF
Pw5l���'E�w�2WW���r3m,OQז�y��9}��7؞y���I^�|���8k�i6����d#���5�*�M�ɢ*�>���뗤�����^7bqRX��+��%��������5NB��Jm�*`�O��o>z�E��iGd�l��U���q�1�X�Dһ�l�ܹ��t-��D�7�̛t:n�&L���>+�ll�ݕ��^�N�s�Fh)���6	���U���䠓�J�-R�k�(�S]�	/�+J@ܱ1$���Y�(�} ��q������l�h��Uz<����D�	�b�7�^v��T��H��&*�3�
Χ�1� �<�O�%a<LM� #�n�K
%aY*��� ���K�ت��
�<�=���;�mY!�j�!rĤY�
�3���������v����o�wa�탖\^S=��B^���
����Q��?h���f�n���a4	ʛ�K���٥@�<����M{���Wù��Q�Fj�>�m��ԏh��ö����4`��T)�0LgX�ߘ��sk�~W���X����`#�(h��w��^}�m�Vm�5���I����7�'w�;���a����o���ҦH:�N�E�b˾v�)\� m �5���s�g充��PKx�+ѳ=f�W;Ǡ^0 ��Z"P���zh3�`�Y?l#���ĊrS,W+#�5H���جE*S��P�쭴�2t�<nh1��Z!@�jVql��֑^�?\VT�ҕp�3���^�<�V�	4�8�71�V�+���c@|��F˃�F�Zǭg����D�X�e	��p+`{��=!6�^�R��ے�Fsy44k_��{Hڍ�_���1�e[��m�b*6���'�ch�=8�����mƋMQ��f)'gfWa����~�Yp�-�8����>/�֙�R@�߃�w٦,#Sn�}F������guWK�R�ZY��R�}}��Q�)V�}�n!u�嬄�H�i��W+�Z�,��q}s���X�Y�	~��>������%�S�>D�����'��3�z2c=�ޯW5dT�����%�B\{�X%�)
7����O���h�Z�'�:h���7H���_g=m؆�[���0�5_�~�7��2b��4����`��>�B6��*_%�T�����m����0��٦�3fb��.76�$�@�_YW3���pE`��[��p*D�?��m�;W�϶Fgk��� �y�v��������"
`~������7��� `H�t9B�Mk;��%�=-�I��t�]�Q}H����S�oz�6�d�s��`X$W��4��ρ�F�(0~���Z���T�c���7ɶڪ��B��N�p܋�Z�����]I�zւ m��o*4�'��w��-����L$I�!&S?��8�-�$�����V��OPٶ�a��Эl�I� UL,�$U*2nD�>L<�&�c�V�1Z�(��L����&(��ɫ�4�Fk2�\,�&U��x���TIc�č�@d���ξ�h�nnԧ��BqӺ�D�w�JMT��ͫ�?�����LE-D}�0R�S
�ɱ�l8I�����#2��#!�_�l'Do�?��-���"yz�D@��X����D��5j�ucMF��n��
j���FS
�q�ߩ�s��v��������	er��L��L�'�_n'L�y�X�N�����}��9T*�K�ͼQ4v�_P����W�[¤%M���d��@��O������w�0e����0�4)�d-~2;�H��Ҏx�ў�����=/YnOw��\�.uv9^	bӮ��mG���H�O{哵�B^�V(m#㋝`�Qqa��Ɯu�]A �zw�V�a���p���=�[�����@��5�$/�Q�4.���X�'.��������y�/e���`_(�����1B.����ʋt�A�p�Z�v��� �r̽���n��7�=-��].n��"y0ix��~���yP��\��k�=�8
�mm����C�@����KA��a]<�H�c8�L�����}�D���{&:c��x�P�������|#� ��hu�M��� ��ɷ��N3��t�E��Xu��Ww&�0�"��&��#i(�����<M�\��vi�F�
�^�<L��@Ss��T���K�p��|�}̭&7�O,����I���$l����f%!��~�0l�b�T�i��7��q�� 8׃&�S#)D6����g����Ѩ�B�I-��:GN��8km���GU��K}�ǻ~'\Y�C�c�Q�+�cg����+4�v����4��R�W��e��z1�{ff~q��|�抧A|�NY���	e/�oA��'���l�����ŦE��IV,�vHe�d��� g/�5jn`L
rab/!ɓG�������'EkT��Ft"���;sh%N��1�a.�f�C�W�9�41�I�1C����#H��K3tM��� qdj>85�0҇��@�$qW��}º\>�?��eZ9G1t�(����ϴ� �e��R'6g��}�	�62��d�z^Tv6;�!K!�դ�F�%E�x����V[\��J���u��^�̧���`ǋ�S�sE�XߌΫnYsw��jmnV	F��@��fO��������[ݒv<��T靕�$���b�D��N�T���W,`۶QPK��.���&�j��2RLB/��X"��P��Ƽ1��&���w2�Z��,�X�#�6�SAΔ�Z�0�[H2;������[���.�U2�i��:>��x�ث�G"�A��ң���b?���j�:��q�(��0�sŮ��*h�2��s�ɔL�+ۙ��� ��8�F��F��x�F�� �U��O�u�jUc�>��Q�֣�ݺ�Պ�t���j;�x���	%����6Yf,��F����A���`���R)�.�y��I�v7�������J�(w��Z5D��i�bP~اA��
���?�::����#Y�ݰt�2kY�P&��z��z�C���/���.��HӁHu�9��|��+T	�Q�(^�d�f���0GcņR�8��:�K߿�DӁ�!	ue��$�u�n�T?�x+'�4���=��^�y9��&�IlK%��hN�l�'q/�3d��d��D��W����3�~Y��3��۶eT���Ƶs�~�9�:����^�0 ��l���>�c��]�Ϗ�vE-��U_�#U��M�"����7�l�,�T������q�剤	�e�<�o
�BE�;� ��Pjx��R�����"�{�w+4N̕�O�GRZ��J�:5A!�A���6b/�p&�8�$�P����ff�Ҹk���yo8	R��M~�%P���~\��V?��w�HRE��QnmA��%��3��>��XE(��/L3����a|B^������Rc]��Lr�3��b����H{���L�q�qw̝ʲU>&',`�Yl)�����.%^�w���_�����,��HEO���NKҷ��Y������C,�l�� �;qS���DKs�`�A/�L�=n�_���\e�Z g�qHQ{�r���J�ܩЌfLa�+��<U�;����xOӗ2*�7����9���n:�>Зj�i��/�~���v.��2�-f���O��O����*��`.�ƅ�)�_�MiU�C1��a��xCԒC^�m%�5��#��5T=�j�:��R�E�W�+���^��3�b������Y�]yq;�*v	�L2�R��v|[���؟���
�e;�{.��*��7S�_b�T��As�C7]���l���	�O��܆;į�X���k�*����ԙ,Ө�-fICߋ�P[�ȝH�py|43��V5e�o�uo����al►�!��K܏��l���G�HW��BaLɅ42@��$px f�����#^��<�C���e�
�8��QyU��>�H�AS�]ǰN�}nQ*��q�|�f�b�>��0�������-�!��/+r�L~e�F,po�,�$Z�Zh��3��M�v�x��K,�if}�՝�R���w�2���ebcw�>�Rz��28B�X	ay��6��/�p��t�Y3(E�+k¶{�Ɂ���;K�
}�:s�#oF�}o���|��t{\`�����DI��*[�>��K߾��㪉��H�f��~�#����o�\������
;9��+Bi�I�`�p����]r��N�aK����l�}�+����I�V7L���s�?��|ٰi���G-�E%i���a
����������P�2<mB<�:	a�����<�r�f�˻���s�!�so]�X�ݫ˱7���#&	/�l.AS�6�NA�u{�h0��T^���e��������{\��!i͸k�l=�e�z_z�$��"BA{����B�e��|".�T���x�^�Zrܱ��d{����p9Q���G���&��wb������B8>ӶzkhJ��8�P)�	Y��sC���*D��/�F�+C���@Q������ʐ�t��/��
��I~���*�N�ﻳcx#� �,T=dK� O�q���,�bfP���G���_�ܓ�� J�k1�؟��:�y��d������h��k��Q|�~����o�P\�v��u`S����$�"7m�2�4��j�f�8H�
iG�_���w���̡��^)4��Xg(�8n`X�H����qlW�[r@�P V(�_;W���&��ò�h^��<yt�\�����>6�H���=D�k�x�C��3�h7�q�^�\-&[�\�Ԏa�
P���up�����.KD�Z�N��Ğ�5����������Xg�Z0����]!���G�a�mB���Ū�;`�:��)���\U�O�m�X�K�mRl{��q���2���n-�V�5FJ&7�P��z�H#%_"����r	��Ʌ�@�����HtD`�Y�8�MD�W�1�scK�"�OӦZ?J[$��kP@$�^'�}?T����fI�AܤP��7����T����0��y����7+�x
�k����"���� �<x��DݼU  >|؊A�r�uyu��f��8�,�w���'�xyu�{"��T�:���F�T�|;��%�$u��l��T�?����J7�8>�ת��&�k�Jmf.MU+�fa �ڏ�Ղ��km���MVA�b5�닾���v7��'�O&j� %�&��ɥc%�Fhj=5Sm��Y !����t�n�"k�[&ڝnw�Q�L@�NNFڳ�n��8v��1�kE��`x��0��*�P>Yg�M�EL~;X���c�Y9����F�fXk��ѷ�;L�V>��9��� ��7���g:j��p�A���mQ�y�F��ȟ����C�(�k���`׉iG葉fY���8�ƹ��d0�HC����eݪz��GS��BD�C�k�-��H�O�nUv�G}\�-�ӓB��<�Q�7��8Z	�\�M��1�w��tn���%�0p�í��L�=_�|�"J=�]���0�r2���"���ȖG�� em�G�����,9#ے��ӂ�orr=�A��j9P�4"��RB�s�Q�O_י�����x+��~��h����i�a�=��/��e"s��xl f����}I��so�ڽ����줖�wҺi�`s�-�xY���-���v����K�Z������ �V��b�g�민�łk��T���E��M9	�n�C`ؔy�~8����������F�=�o��T��'��D��N�Q<*"�=!z�RsKOk�z
יg3��>{MҀ���9�=kZ7���Y�,�\(�S̃����l`L�7\�W��?�a��"T'��=��3<��́P��(QR�0�m.����`�VT�������x2VEo���5m>j�Idi7J6$�/~c<7PX:����S�Y�T�{`������3L�Qq�>��ڵ@Wѯ"���^Z��a�J��'he�澛|j�����ܽ.��]���X�
�H�2�_��jp&;����e�-�;<�^ҽq�TWt�2��c(�R��	��y�V�hzl���Vw������]���ؒC9B��G���������}딿[����k2�ӾNH�H�RHs��\���f�@*�$�� �-)g�G��)���b�-��6��Sx������4��z�|!R�����=v�*�m9�k�?�z�O��[�nv�P�il�SK���벑�OE�U'�B���bx����b�{�Ɵ�rg���(�OI���3��l���!��$W�C{U �k��&A!:!8�T]lVy����)���V����(nq*�Y�҈�[)��%�m_��=bb��U B-��m��>���`\f��7<i7ll;$ڕ���_�Eb���+	.�q>3zQݝSS!�8,+}��m���S{ʛ<E���N�l2_�g��Rø=��]l�$6d���곕�|F����0Ͼ���a�JPa��R�J|G��Lj'\*�ّg��?�����`�i�s�*>f�0���,�#'�AS0�a\�hJ���N��F�T(u�"����h  P]�i�&���uQ�&+A�M�].f�0��>F�� �����޽+����|w<������3��g���=�c���v����kd�!C�,�s�)I���;fW%�}�=ݶ J((����̡�m��E<��Q����P���Ӿ�������k��;��X�j��q�L{.�"�B�A?6E�I;�E~�jZ��;���������!&N"k����}��D�v�xz��6�s�i&A#E\m��-��m��lǘ���_���#�^甶��P���;R��gĶ̽k	Am�!tY�jh��Ρ�Y;�B����	�����-�J�M,�hG�C�*^��/0m*{���ބ��x)G�� ��JU�i�O�Zȹ} �-�Pu�1}�� �QT������dY!3@n�u�S�S��9�-����|�QΆ�%*��������o*���<�*:�bw�MFk���,�"�8��/'e�Pd�^���bOB��%wD!�D>3[b�a�� �P�j�'��(��]�8�Q'Rp=�$���:fҹ��7�zD$���p?^庠�"4r�����+�g�����5	�j��u��sq�l�{��=|�+�(Q�`��f��l��Z����ғ���.���2�nKF��Q*����ݾ�K���� d���ۼ��/Xc��}�I�[���809{���IVG*����p�r���=1����[��A���}��/�em�E���5O��Z�e���,.�|��V�>w���s[�9;��0َ~sJcI�W#�t�b�p�0^$��P�v2�'�h����-ԙ�!$�,t=��	���{/"W�d�v¼�-�&��U1�h��2�~�1��HeRi�)�5�(�I��`lW�J�A,!`eia�gPːΪ������p� #�8�
6WP�*�#i���ްh0��!�e3��t�clrb}�ɩې>gm�|Ox�w�bP��Vڨ�>k����z�}��Li�'n���i"��s���ȗ���dA���@��IM����o|�_��H|�>��~/@�]�K�$r�TI��F�C>�*���~5�GÌs�u0\2�x(�򰪨z�%7��>���{��m٠�'��~}�h4�Gc�p͛�ٱx+��cS@H�{�5����a�����j��Wl\3����J��W�4�4ƾt�6ewZ�z��{��'4�x��tK[c�e������(��ډ�Hſ]# �G�z��ߩ)O䞔���[D�
TU�(�a�h���W"?3���_j�t4RNZmF�:æ�k��d^�/��97P}��)��7I܏�	�~�睍N�-�vW�3&�)l��k�R�� ���LH��&��
�󶆰$R����k����r�@���y���ْ��3��@3Q�Ed��{�cF�N���W�ˤ�CEӵe�V �Īae��,n��v^e-��7�,=�4�/Z;�)�tKy��Vu���Ê@7b�|̘϶��$lC�|������9/"`�pƻ��~Ꝕ��g��b���|8��V40~�-��o�j��qY�b�6��I9�Yc#Y��#�@�Ӕ�������4|P�'a�`�p+�t�is�qZ=!��
�m=g�(V������r���Όq�_��g�Tz���w���|D��L|p(�}�/"��Ca�I��~��V��*}��;��2�Y���Kh��F&��0bs.��%��g��$u�E=HY��	�pp�H����3��~w:} �)_��Z0�
%+&B�
�q_�������}ًl���Rcx�e�d�^\$���5� ���F��	p� ��E'Ʉw�5���3��`�*�٣�pf�v]��A�	�:D�4!b�����A������W�t�lq����R��	�s��M��=^�wDN�� ����\,/�L�YH�-�V��C����㯗�t���A�"M���6�,��$��A@[�}�`��~�ş�V��5�Bx��]ړ��y�w_��1.3E�R���������:�X+2�EUǃ�ͺ�/݆�|�2��KH,�)p�&�~[��9��e>��ɘN̪"�9dG���U������b�qY~�Y�d�ҫ<��_H�'�V���z����x=�WѾI��-{�k�X��;�~�%��)�ł�[�8Z���"�W�-��� �����X�D��e�����[�[t�sY��*E�'DR���u��h�Dv�-����k�2:wə'���*3������c1d��"�7�bw'\��?+����fP��Ͻ�d{��ۍA`0.Q��8nw02���:�@���DY�y�ٳZ�����;'��4E@�X��s��Ji����,�F/�D:�em?��"/��8z�Cdn�QQa��6�ShHG�����`v�=jo�j��h�图�VS��~�+y828�d�L$4#C��e��+��x� tCc�?}��H������k%z�%��]�|cɧ4��L��ta��ԪyW0�em����A
�ęe:�=^����\-N����&�X�Mp�+��Ks�����ϋ���Q̿W�:/��C�؛�ժNޞΊ6%�sBt�u�;4�NJI�^m�(�����V����k�W:=�F��{��LY�;���7\GF$�3'��㝈�\�!�b0܊�#��Rd�h�<K�^c��$�����u������q%������X[�v;�`W�@e��:a��\�w;��ù$x�����~P*^��<����D�N�[s�QH6i=�r5��OK�|OMsu0؝,KꚯA876I�,{Ǣ����k�*6�2W	�J<��As�W�'A�H�π�1өP��3U�!��˶'W莳-���m>�zj����e�s���ݟ@��b��Ҏ�Ë/Z�-"�!�&_On
�%���WM��н��}�^Wb��=
E�e�B��p;�*�5���F��������~�qɔ:�G>�O��A�cwc/=�Lc�՗K���Vω� n��Lr�>ӟj� ���3d�	p^��{�%�pұ�b~���'��5���}]��bΎM�Yd�iP��J@�0u��#�+W)��
�sa��T��v��Q��T��d��5#�1�����{�x�_7-�O���	�h���{k���	�e@3�J����RL�稊1wT�</o���7m�T��T��!m-b=6:!�p��|ū�$9+�m�T(�	��_m�L�N��l��)@�C]����5��БTܱ�b�����>mt�vO��˼�L+i�� :I[���!�D�Bso���������byr�W�Gj�:An]�m��D����s�N�r��#FpE�ɜ$�D{S�Ó��C
w&��,qoݱ鷆�uf�(X����?JN7I)��^t��̴Jp�&-E.٪w�ʌ�-X!V&Xmo�RK�!�m.yR?�� �9�'~"�_��������hu��`ߑ*����7y�'/�@~�Ō�_�_��l����W/��$*��t�1Qn1�уi�d?��]h�Y��{�bE.���A��w�^��榁h��]O<�B��a�� lq�$˼0	�3g����\[��Ǥ	x��Kj �Z�x�I�^�F�`��ktLf�`�0�	��vl��� �}��|qV�o-���J���DW,�6�Qf�@��ڍ.����K�*\ ��떿�R>�+\n�Wȼ�$}x0�$u���U�䪜 VMX����[O�0��X|v�C*w����Y�V;6��a��ÆX3�\֙���ޮ�{���q�����nNpZnw��N��]��OU��m�VF��xBd�52����R�a�i ��j`D�hCZO���(�$5��p�Y�}��X�A�s�d,]wd)�zE('��N�M1�<���X^6aV���Ȩ�>K����jN��u I�[G���{��:���[^��죲�V<���nƏj%�[�	��E��,����4�B����ю�`m�`�7�:t��f/�L��PA�<�!���#���D�+��qإ��^����=́�ñ�^M�v'~�{��v\�������vg:��$�|'�"�J�w4�D�����˘FAM�������3lp�o�#��ۤ�g�C��8hU��	����V.M����8:���tqUBt(nW�?)oYF��$��?n�c��0�L�_n�H���vn'�{�����m�����qN��a0���Ԅ���W�֮]����x�~q���P�ףm�X����������<�����SF_�F�D'9�����=��}�٤8f�	��or�� S)a�^F�~y�X������"Zn����Lg���I_jC�#�BP��3��(�V��[�Wc؜�� �F���Ș+�T�r<:j}-]�����Gn���,K��0q��,&^�'�#���?�v�m���<ι���s�}��X����hwH��?��#?j�Z��ufT1�V4f��§�
�����%3���\󵣗����JX	K��U��
K^R�|��a[M1�#�Y�8�H����J���7��$���)J�ȓ���j����2s�2���;�E�n��IDg�@���>�Ǩ� ����4 ������?�8N��w�0�b78!�����ƢN���g��d�~��1 kt��	sX����߾����|�U-T`��Ŵj��h�����4ڤȰc���%�����K:%�>��+F�d��r��~X�g Jh��Q3B�<ׁ��/R���]�Z�7&#��\\����{K�O�ՔdPh"�|_т��;"_����;�|���}��3�y0	.͙����T�����\�
O�iJ����hB�E/��&:�z7g�pۛ�: @�DeRlKĸ�n徊3w*�W�|7K��6>�e�3���!֔��J"J
�%�]��W+[B[N�DlT����_�i�~���lR~o�lA��G�K��աl=&,(l��Y �����ҟ?�M���P1&�M����q�[���R��LEs��ч�r�4��陳���٩å�}���C��{ǯ�/�f���$KX�S�(����;XyL)*����5��D[�S���$��lϿ���5�\���KG�a,�������&%�����U9��q1D5&�@+��\P��כ��4������{��X�a��\�Ƴv�J�r&Ӗ�@�4N5<���/���p ��<l�2P;) ic��G�0M|?s����@m �uc��J����������u'����8�d!3` >L�g�q���4�lu�@�m�����O�J&��5F���DL�L]�]z�� }I ���7(@@�<n��W�N={�-@C@G���7��UC;�F��z9k��ca\��;՛�����s���xU�K�R��gQ�X,>����� �Z�����p�������[��J&`d|z4��=W<���(����ԦȒ��ۏ�"+�WP����Уf��������<?S�U��0����H�������oą���wR�f�q�;X�,��9�k�ڈ��QO��)j�r,��VdV����H	�_m��>-�W%K{�b��[�W�R��,r�暯�IQ�7�y��X�[��Z�jW�[�n2 |��y�n��:@H�xJ�����߀�?y4��l�ŇG���Į�BY+�S�	���?�t$�u���"�ji�̞�Z�M�H.��f��c6>e&Urd�)��J��w� _M�Y�y��c�hӱv`X�g �Y�3R�ODDx�D��D*צ�U�}���Au]�˩��[��7*��δ��Y��؄%��K�ɞ&(� �2��П#(����^�3T��{܃Ci�G�l����EL�qV?I�r!~��7�w)5X=ͺ�_���)�a���n-vf�e`/5��V�pg4h��{5������y�ث�se���e$%���/��[�vyx?�\A�z���?	{��[ӵT�ґ�)�ي��g��1�2�k���+�s��A(,�2�{*;M@�1����n0"4Ǌs��>���ۿgI9`x���ge.�ǹ�9<��EL�4�o2�y�9��U$��(w�m�X�hd7i��nĊ��HG�~D~3��~�&�����q�?wd�n&)��|�����E��O_������N��$���%�g��9�s\�b��o�`k����<�Yt���U�,�Qu�,���fC�'&��nL��H���Ye�w
�*��h	�����#}:iGO��zJ�V}���y�{P}�>I�O�R�8�K�K�L6��"�L�RM�%��&~�Γ(���O�`�VQn~���u~Y��(�a���C��r=���~�MbC�P�Ql<�pW����1ꅋ}n�`��@�k)�b|gk��t���@R^�x�_G�΋!	?K��u���@����
��i�t����b�
.� q�M���H_/�^{%��%�KD�{g�G]��0r��3	*� _o���U2�ފ�Q������NM���E`dp=Kb \����{Ъ_a`���RN�#(~ǟ0�d�8ࢅl ^4��I}<BP{/����	���M%����`�{�\�G��.�{l��-[Hc����D8у.6oe�WN��}�q��ӕ���O���<K�34�Q�t5lV+_�HF�g?'J��)�N};��^��r#�T��3_].&ƪ�1�9�d	@cg����s�fe��J��7�|xćg�B���[�Q�ҔG�x�L3& ,��`�F��f�ve�oh��� /���9ЈO��x« ��>lTQ��Ɯ��wl��`I��(��H�����̋0�Y�p�I�=��M�E�d"��?�����x��L
՛�0�_i��`�ļ �8��(�\h!���n���1U�tȣ���������x�m��L�.���s� �wӟc�� sgT��R�8v~������$���j�4�ʤ�jB�&I�&��Ү���]T��f�22�0s�`��ѓw��)�\�����__�[gu��,����9�ʑ�G��R�@��q�T�L�)P3&S�Cw��v�0����\���Ҋ9���|�WH0M�٥�Ԧ�j�������'�A�@�}���+ʲ"E�=ue���v��l���I!��d:
HBѾ����0�A��U�т &ґ��g @����eA+wxn(�b�u���in���O&�V�/����^H��$|��9�3H���P��h���7��N�BJ�%�}ʉ�	�y,�p�Y�=��7��Q!��=��I��Q�箴BBFf+O�hu����.O���u:NZ�q����ǽ��[,��Gi�f��V��X��:�9>V�B�{~e	��%R� �IgH�o��GY�LCq��op����s���g\��E?.B�V�0��R�b��X�)�؉��m9�_��2�[֘�Bf���=X�sb�����~�<��Ng�O��D���%�ܤ��}0ZtBE0�K�s��h�������*�r�
@~��d5�=��ԛ�.S�z�'��X����ۻ��K-`Ч"�5�0��X�����a������l6������*C��߉[>7B��8��t��yu�� ���+]�i�n��l%sf�Q�aQ�L���ԉ̊7Q]��������0`�x��2 �'�ƀ���Ϸi��E�����8!�@�Ҝ����\�`yupl�sT�u.+R�~�GxY���*@o�~��¡q]�^�&�a�悟,�7�ʽ4ҩ|�{�k)r!8�������W��&��~	�T��/=�/D����|�R�p׬Q/
��m����^�� Y�N���P��u��z�N�gl%�΍�o�[�|���du9ш�8�~�|d�xiT?an�=tE�Gv���)��{�G��y�'�Bb �o������1ͻ�>��+�45���X�uش��C�J#�&/I엄��9�4~�M�D������t+� ��J�]��i
�]��'�c��ŎǗ��� �T�v�eG�@�j���C;S�h�KZ���5e�f�b��P�
o���*�iz�X�! �j˚r/D
`���K�@�����m�7!΃�F�� �%w��yՀ03�@�u�`9��?gd�M�6�V���9������4�}s1O� Ԙ{S��#
_�rṯ��^2�_�t�I�0��U��N������(�i�����9�"��_術�ܶZ���U���ؾ�T;q��_��;wm���i:��r��ڣ�X�/�;��aO�]8y������o��fn��Y͓h$
�w��,gƸ��S�$�K�Q��A7��S�#p��uco��]�/�=o�����?��$��z���YJ��-�5�d��L�3o���݉^aYp���8=Y�J�¿K�'��SzJ�Ӭ]#)tc�7���e���\�c�������1K}��h���O�|��c[��ZD�'��@9`H��f� ��a��K𵑬��a��&Ft����J���|�	fӔ����'-?�*���j;>�U-)�IBP!X7�������?8��]��"��^KtBC8i�vŶ��;�`!h��f�)�#�8֖����[�WX���äV����I������`�hn"�J�� �*Q����',��6Z�����g�Ŧ)� X��"�A1��Ϲ�|���qw���`P��9��qEEB�޴�c��L��B��H����҈!?DA��yB͹�jz��1�m�1��7:2J�l�gD�a��0"*�-WA��V9��v�s�������\3&�O-�@_�G�Zx�V��鯝C"������n�V�F�e~yYnr�8S�\�c��^ii� �͋�*���(c�!��:n�������_n!GF9�k��vzу>��4��ӟ�gMN��'m)�lQ`|>��������u	���P�+�$g��?��U_�6E��D
�@$/�n��\�mx�����]n��zH��N_�<cRe��b4=m��Ǩ#sH_헽rx��qF��|�.z���\�(4�(]���H�
= 
�Ƿ�֮�&p��ܥHBH��'�@Q�$����X=��CS�"I#d��0�>u�d��n���lQ��	o�� "�R��# �ɓ(A�,U��	���h�io���Z�����3��������U\��e5�(�z�Q*[y�����2|�V>w��8�p��p�|��������3�u���ݾ�G��;�a�Uگ��_@ͩ�2�h�I���~��������kx|�ܮ��:�%[��ɤAoУ(�M%�6nm�G�VR�:���We_��-϶���@@���if=Q�7���@�<K�
R���s\�M�~%�nG��&�I�e˿�y���7 ۈ[����Ѻ�����sD{��UN��I��l�|�/�m���b�������j_�q�
^���֜R�{v���r�m�ҽ��T��6�#nH����tfx�8���z|�Bv�L 	U�-ϫ�4B����^	��ʓ8~*��}y�Yl}�Heh���k~5�"��u����>����wUV�L�4�1�����k�]zp3��d4rh���GwtVw`H����Ä�OY��t�������Z9����4G$��ؽ�I3H�U� ���b?:s8��RVwA�(ϏӲ�e�h��a�D��<���WFk<īg�k�f"����=ek�D�_c���i�ŤG�9GQb�I�cS�-J�K�M�?(�j:�Χ��4S}��}���X��5�!;n��a��㽳�?�vF��iT
�x�3��ܷ@�8~Kv���Oe(7.�otR�c��̾����mei��.֊��l�֠~!��`C��R������9T��Hč�U�]��%l��?�5I�2�L1_��b�Z':t�t�-�o�KXU�#Zр'�9Ǿ<����S��T�L!�?~�;��!Hj@a��>�a5_S�,�怟Ы���)�I�%U�8 �[|��vI-R�`,ږ�EN��Yd��vB#�Z�rG���h�)x���M�
���ɹ}��������<t�����ev>|̔w���SN�}Vl�������-��<���l���Ҭ�%��f^�?���	�D\?�!㑦卣���n���ݒ�d�b].;_��o�\v��	3��g�ꌀ#��u)��HKE'�[EwYg{;k��-<�(e< ���
�n$n]���H{��CJZwb%U��{�,�$B��9o�[����HM��R�A�=���'��-��8�˴�����Bx�8[�;S�`#jvS�o�{�pc�_�P��/��
�GA��QCr�O��.!�R �e��^+2'�u�� |D�Z`�4��	�&;�Уl��}�]�~���f�'�s��u�� w��� �OV�?"�)��q��Y�C:8O`����Z�6����[Do����$Nʳl��J�}���yF?�w������U5H�i�Ю2��؃2١�f_r��Wᘌ1�pde	6`YL�K���.�<���J�+P0M�U<��E?v� ̎���O��F��0�2���w���ϐm��b*y�h�0�k;>Mi���|h��ִ:�ډ-3Y]g4D�ϳ\j��c�T����c&����]�4k�/f�tz�+��� ��<I�@��v9b��}*(q�E�Ҥ�KY$�7�Ĥ�vAE�&g�ն�$U���B��`��
�mH�j�C��^}��ZzX8�+��K4 5=�w�l�PM-�99�*�9�[Ca�z���m�iK���x�G�4=��w13ʦ��V��<�f�� ����<&^�D�`��;����.�)�f��1�^sr��U�~�:�Sak/�"��=	�nxosߴ���XU^�dlœ**���7@Igisr~Z��W���u`#�ܟ{n�8霁�,/�)4v���Z��8ד6�(1���ƾ̵ޏ=�X�l�6��o����q���0
4������x3h�:��!$������}� Atx�^�j���@Z`XN�,��W�,�i������ԙQJ�Q����9|����>ō�F����V��m�EX�ph��4CfR�^9���QO�} ��[�%�2NJ��H���;Gz<����}ٟC���]Ey�Dܶ;`�#��:#�d|�(
|8Z2���x��E��OZ�ֲnG�Bu�m��'�b���m3�¸YD!ԕ<K�*��g�����[!�	��Vߙ@HA�]7�:SL�;,;���$�d��跿�7�NGMB�}�<�� ��I�VR@���$2\|[aLn�+I��@���E�읥He�NP�u˳����w�:"NR����}�R��,e &&�g�s��a�P��������ܸ�K���=<$}~p��'jbhV��d<�r8�ɮ!(_i�F����j��)q��/����)6yY�[*��[Γ`[�6oH�d2��by���)�^��g����GAv��%�
I�l�#L/����svV�.`���0��+s,uD���� f�
�`�����8ٿ��akK-[q�h�><�U�N�N�*�� T.�_��Z�r��\)�ea	�]ųg"}}]��<*��ߖ
�%���J�0��ȗ\7f.�� g	A�!�g����E��L���0�&s��f��wi���%v}aN)&J�YеזaF*X������ ܣ��r��.�s�-����uQͻ)��/�,�-��m��Y,�qڀs�+�7�oO6D׸��FO�[��ڥ�q<Eg���!e�w��a����+�z���3����"��uA��7͠})���OHŜ�O����1c��~{����!s	Y���Hů��«��MJ��SS$��x�Gʌe+v��YƷ/�v��R;����3�*�����X��1�9�t���pD��D��<�}�c��ri�Cȩ��aC�-�Q��J���[����,c}�"�.n��`�N��k�T��d��km��f��M;���
2�a�a�����T�o��a��~�S���}0��U�F{Od�:��$VQ\�!MZb(�=&�L����ёd�/�=G�M$�l��l��z����U)��dx����kĐ� �*����E�$�_�D@�nL�혰�[
S�BD�#���Y�R�uv�d2��A���� B�赵���T��$���pm��/a�CеXٌ�$^aI��|���YI(�D��9������:xU'��F��	�Ií R��x�*9������u��sE��aamǲ �c����ҫtOp�%���߲�.�;�Fgq�L��k��\^̦O'5V��}��ID�m���-��Lr�7��'�&k}�QJo@�6y��ž�k��:�.��7�'��}s8W~b�%�)��sǮ.ѹS������L��D`R1��j4eP���K�t�����d�=�x�s���V�̝<��Եi����'���}�;`뉖g	�F�;���I�,��m�a2�bk�� ,����:ǣ�Q���F4_����b�e��Ρ�:2�%�j����i�$V��Od4g#[%��g&��������U��t��o��ؙMw�A�;�qƝ+$�<z��}#��hb�lv�MĘ���iĩ@����̀%V]\ε6�+&k��()k�f/+��0�w��%d
��1.����? .3��C��]�Ԅ���d�ǄH�+��Ka�[(k����׀�:p�e��`m��0j���4��W�N�2>YVT0W��T������ �N�F��a�
��-S�o�FA���	�7t��{�C��ϵ2�@���T�A�$U��	8e?1�J�S8$��L��p�~�E薟-g����th�T�r��Q��l��T\l����Z��/1�����R����!f�6_U���Gԃ'�aJ6�������ko��R��oق��G����r��R��8��$h\
Ҿ�,2\}�C0��'b4��Z&v�uh�}���^�M�$������~A�<�>�S�tv�N�7j A�Rn>��O�`o�dF���J��E4U�e	��Z�w�il�1���\��o�|,�x�g�i0��v�#�}D��^��^��!�Y$`p��rP��4;�R�-�X�X�������W$$�����``��A"s����;�M��L�z���5�*Ѩ��	7�R������d��r�Ҡ�����7�%���ƚD�O#У�J�/�}����3�NM^�E�m���^��e���؋�^�q(Ubk(L˺���$�Uo) �و�mG�_�`�M����7<RE�c�Q�NͰ���2���%m�M�	����F�b|�#�-aۅ�s&N��/�7�k�3�8�.�r!Ǌ}�쾞sxa����Gw���j�������CI��R�Rt��x��4ee���KP�$��{b�3��yV��M�Nt��	�%NE\�)џ߽�b{�g�)6�2��^����d��*���/���Qf��D�MуIg�â�>���ca�o���GR�c/���(�8�V^�#�3��B�C��`��:�v��;��E����0_��ܙ<Ƣ��
�V�D��4`zॣ���o��X����$"7XrK��(ʯp�3Sr����a2���m�h�L&?���߲���O}�ׯ(����dh�c
��)�v��ǆ+v��|21�)�R�KI8��o���c��'�	�Eg4�z_[�d�~>��vM���x��-�^�ENV���n�Ķ)���%� �d�G��	�|[����*(z��)�e�(t�D�%d�bI�
�k��fs��I��$����*E�o�>��)%c:��mX��!�q��ä�36+�;�e�;��Da���x,���Fv�44�:��}g�<�ܻrץ�P:�j��H�lIǤ	��gL�`�.B��)JU�t��w�7h6^ r#w�3�챊�'�x2��	��%'�W�>$��4�l�O�M�~=7I�,H#M.�3��N�I����Jm�0�t�{���Ec�N']]�y�?3p�mW�A*z	g���ȇ��b
^���O����S�M��DM���y@2=/���HB'�4�������߇�PWE'�S��g�|�5�˰2��s���$���戡�a:��V@FY�ګ�z1��v���E�pѐ�A��Щ |l�ti����n�dJC��.⵷s�
�e�%�[3�x�r��(Vjg�Kth��}�1G�W2��K֔4[��^ú�ޅ�s�/����)�ʕ+e�[:+�mZ=�g����yw'2��)��I������u�Q���k�	��(�"l��(�0]
Ks�Dec�$R�lهIg�9����3�oƧ��μ��7��o��)�V&�Ci�ho	4|�Rd23v�m?��"H��kf� .�ۤ�R���X�����+TL��!�+�ї�ާ�4F��V���'��Rc�M�'�_l ���ִ�l��@��ȱM�1�j>-nA��?���FTϘ���C��{Az��-�.��EҨ)K�B/j����T0�;��m�լ4����?��f�.��~Ⱦ[-�N�ξlrM%CV�D�E?z��l�
���b*?�:�ُ9-��u[~.��ꦌmnޔ�
QM���(����D�j��"@5u�i��q��v1� J��;$��Hz[�s��wC:���#<ګR�Sh��m�/�x����%۬S�~�6v�zmh��t/{Onn�p/%�D"v�nE�h��.��9��.11�3Д�
9�(���ϴ=H���ѥ%���:���c_���wsbH�z�q�f�z�ɞf��/��'6L��A���`V#N���ս.�h��U#8��N:|���1�~�����]��q�D�K��A�x2G�����G�-)���n��b#+������)�[c��j�2'��=��u$�4W��]5%�r��o��u�r �7`��U�o�J�e��V�z�'G��m<a��yЎ��#NR�h��0�CY�m��\�Xl\/�@J\�+��e
.۞��UL�e�bI��4�]�g%+�hDm��7Wt��u	[�7�ȓ�Ъ�B�X47e�.�aiׄ's����_K�9wr8~���,�zm�����������m�&/��σ9�r[���)pLR�~�ozo&?y���)d�6z �*����T[�j��:J�6%�B����kи�$N#�v�Fs���<�y%
���U��K��ĳ���У���pʀ�@my]�bD�+Y�ўT�����>�Y:ں�3�\i�r10}g:�%�6�䜓V�䒣{G���ZK��PW|(*�*��	p�t��l���j)�X?iY��l���V!+Uߌ��8-E0M���_�բ >c$ipJ	U����Ƌp9�ހ�#��نG�0�)�R&�i�i�����R-̂Y��� ��-ocXAN�)S")S�g�=�F��K4O���	'ⱹW,?�xs��Sr�m*l��F�垴u�%Tgo�D���<�áJnK�����<v����a�s��`�����MǼ�R�� ]��J�{C��+��m��^����!���wT{@6�8`����`��є�<��\�J��u\�C������{�����Fw\(j��0ab ���L��xF2t��]_��uW�!f���+��}��ϊ��@G�.i� y���!��O������ػϔ�6>�У�o���+����J�&�(m��-�"!)MW��uSD��
�[R�H���!���䊓V�a����ޒ6B��n�$��o�3=_�f�J"� �u
��I�j}�kӱMsReg�b�◅]���hJ)� �J�w)R��qT��	hp�#�&����Cf͛	.[-j�������O��
M�#�<�g���?�E[�w3��^/";�6zc��W����%ЎU�ű�rX<����T�&mA
ژD~~��_ٲ��u��"5��м4�{s��JGp�6��:��[�S&v�oV��K�z���5����O�U�2�: ����������hS
�@Kl�w���!�g�^�y#��te���4� :L�Ζ8��c��F��!����F��xg�ۏ�nv�e� �7bA�(!�m��p�Ԣ8��=b��R�
v%�wF�4���sx|s�~+�f#vqt�jяĐ'G$�DҸ�*��u�R�#$%P���4�U��~{N��Yv� �E���p� ���}[-Ν,�^�lĦY6�[L���]=ͪ�������B;�Jt�WEA/"�L@�ld�:W����d4녌�N�:$����Tl��D�Uґ��p�I�:�2U�|�c�&/�a��}F{coֺ���J=>9N��;���囸����r͉�hW9��bP��Z^�@y�u)�}���h��z;*}w�Ǝ����V�����A�(�����oK��p�B��Z�������&.p�:Sy�L��	v��T�¶�M�k��GB�Ģm�?f����G�(�s�MI��-�R��D��H㾯��Aw�o�1�&A�Kv���^h��B��G����z�yh�#�ꕆw�%�������-�&i��Y\�C<��иp��ά�����I���.	����`�����$��4�>nt�(
�&C$�Q4[}7*�Oti��5C������6!�I���f���4d#�����Ng��ivl����\N!v��ӕ��`�l�p;�}�e���q �N(�x帇��?	�G[/�Ie�Ȕs�j��N��e�~P�L�6��52�R�η��J�H[�aOJ.�2&��\$I�|�|q�oܧ9��1�n%c�Y�4,%�~�����'ȀHkm�i.�%&Y�L^�"��C�`�o\0`%��Y樂+�G��=�R�r]��E���#(�F�x�!�]�76��s1�p���TpT����q�J���F��.�?��:����ٕ����N��ݯ��Q����9����N̐֬,+D+�M��y=�i�x���򠥂1ϜJ�WC�⣡������>��Z5=�����C����ik>v��+�]&)"2$d��.�.�X=q�bߏH��H�/�������bEGDFS<%�UTu��'���y[8O���m��/��7�#�D�L%��p;�Yζ�^�B���t��|�m`�j�Y���S%(Wasu�gx�<�A�A�y��q��
@'�ⰾp��~�����uS1-�_�$������Y�+d��3+̓��c�ư��	ҤC���d���0�ʹJAF�w��g�!�å�UC�)���sV}��M��嘡U"m�{�]��eل�r��[a�.�����ևWQ8k��Y{��>�ι�4�\Կ1�%��r�S���_�ݼ�L���(�F���%u�YZ)$ ζ��,yŌNq�M.0LY����9���Ͻو���|��"Y~F�:�_���7��S�T�"N��Q> .Z����}���>~�X��N�'��M��{�`��;�r:��VS����[�	�e=�@H�r�=,��%�,ka��7!���N��@����u��0�y4f\}ܒ��Zr_V@��X,�_G\�T�P��F*MO��j��J��RfiL:l���;1qRh��R��f�+�W�0v����_��C��g֮_�ln尕t�]�ڤUo�]m�Ͽ�t �(�a��T��i^��G���=�p��"�y��b�U�t.4��ܰ���V��M�%�2�a���A����|�h��_\�	:���K\�c	�3)��ʹD���ɧֆ��>_LI n��N�}[m-�z�>jeD'y
j���)ʵe���F�5~��K7�N{�n*Q�=��<*�@��'�N���
k��a�����CCu��eC���X�b�x�WB廸Z4ś3/��3L����@QX���� ��lY� ꌱ�c=1��fQ�p�`��%���#0ڈ�;�̻_KNfkE�T��b2\�- �Wk Q���+��C8�P��=�k1��Fǃ�Du�����,(��$p��!E%9dK�N��WG�I/ ���(�4�|�J�t����P6�{>T��7���A��S)�AY�3C�^�U�^}���ߩyM��?i;�j2kY�M�Sc��e�J�|<aV��=��	�e?�6�h��
�A����0�����j+��)����q�P�l��<�G8K�u'�[%q4X����6�-��=�$zU�V���hyw�@M�+�:=�{I��e X� �b|d��#�JKUbPK�Q����ܮ�[������;�~�����nZw�v����; 4�U���[��	�>�.�h��(Z>{���P�e�Ĳ�;���ӹ��F��6S����k�(��w�ߩ7�G�V��ҍ�*�)�'���S݊LT�?�I���|ȍ�����J��j����.��ݱ�-on�%9�5}BXqV�!��;�i�B~�-�� ռsź�J�R�f��!8h�����P�!|��
<JJ�1�����9�&@hN���a��i�vd���ʪ����G/Tg��F٥��m6�`M�:�Ca��=��Ft���<��~�ly$L��n�����F[y�4}��/�1���b_?Pa�v*�a}��x�d�chNPCLF���-8�8��:��4'�sg��UB�����;�5NG7Z^�G�y�yE����E�m���]��=�x�ϱ���cEvG���36�)�[�`�[S�y-��?]�CbG&���ku���RD�H�w�������'��<:��b᱓����ڔ؀^�w©|K�Z�:Q��-�5�F-�0�~MM0�,�ŵ���(x~�Q�L+h�<�=q�Xg;���+��m�`іV�7��щ��^�J8��<I!��
���r�f82o9�?U�@�_�C���V��IV:W*��ji�,w�/�t��s��}��!�uA�EeÊ�	$�Sx"f�x������J���+��n�Tb(2hLV��ʲ?BA�2�0�+���]q�yj��c�^���{,������k5at#�|�[�5w����}.]�F����YvJ`Cȿ@.�.0�||.җ"�*�6}x��v�P	 �-Ֆ�<���*sh`�@�>C!��\�2�@F��@s`����<��p�5�p�J�Uy.�.���v57���p���xG���n��ow��2��r0
��_�q�Η��F�%�~�kG�P��l���D�2�8���rKG*bv���N�g0��6�<C�ĩ�k�0���iC�|��3�*D��_5 s�fB������
ؒ�I,Ĭ���+B�*�I�'l-j���Ԙ��s @-Z	��=�����;xp�]���������4���Þ[�"��^3q6�P������~TE?Fyk�7(M�U۷�tP.c	�I��̲�������V�s��+@b�jnF���=�Df]� �����˩�A+Ew\� �C�l��-�S�/^5;���W�ၜ=\��Vs���rE�BV��P��L��[j���T��/�"T�ꑃ]w�i0����go��ÏH�}�����_[lJ��g�B��}�H�R�r��H|�/�v��?�6F�Oa���@��I��v��+��F��q�*yL�%I��q=`sN�T䬺
���!�7���~���`p�z�Q'��n��Mp|��sF���%Z�K&q�!�%n�l��<nw�:ȤJ�x��/4�*����r���v}j�~(̔�2^���IͷsBA1;$(W4�f�&k����VxK��3��1U������۳y����Ɋc#���qE�����V9	���r����� �vd�E׮qo�����!!�*��El�&��j���S��.�xM/ �X�t�6B� ��P���:Q��0gY����wL���w�9'��\AM�,�;��t�5q蟼5AÈ�Z������5� ѳD�AiQ��g�h��E5�����Ҋ`���>0�#S?��·&���=�?�O.�`�Iuu(�K��S+�{��Ǿ%�6�j��;!B��Ž}7x�$^�8�%�< =4��r�� ���.��/����a�$S�7�A/�X?�#�%>i$��D�u؞!_�O��m�5
�[��r�D�Fv7T6�Dƅ��i�wm����8%��������҇���q�z�X�b0���+RV��@�]����d���f֣.�pC�e{��������ށ���rE��Gjɡ>�ѯy�U&����S�W���<L�`@�%a2���������ѧ."_l���"Fm��7ɹ�5�i=�l�zBB8O߫���#uN{Vh�f�,5��Z��W�
���F� �eC���eN���>����[���ڽ`���J��x�����t+/��+@�;UP�c�&!E�w�S����̅"	�w�9��C����X�x726���Kԛt��l�������p��Ԅ@���2�?���.A�����J�������x\�Tv�÷B�70�)S��G�}Gr���������qb�?�=����m$W\��x��k��'0��"w�Jbj��#X�5�kqv���PDHì|���W��>H��!O�`�!�w[�1�Tݔj��ji{�J`I$,�Pڕ���5��������.�������YE�T���\WJbe�"��B���>$�h8�'d������1zz6}ӝHI���ǝ�Z^���je����I��$�M�h��I^�ܸ,[,��^j5��-dG∶��=02.��U ���i�3BA�"�̬#L 	�zc1���d<j�n���a��O�7'��]��q�'���W�W����Ng�R��F�����P�uD�5 [�<z{��H[��ߝ��} �iU?���5*���9E�r��vNd9��l��ex�����ǫ�����=,�¡���ȍ>���W1�3�}�[�V�ELC�훾G����K�U�m���X��9�s���\aa�@p	 ^"(�+A�^�\���dc`򌶪O�`:��V�A�����!w'$R�2c;�lv}�E�w/����y(˘��;�����E�-��b�������m������`�a�")�Iu?B���P�˧���m=z}�E >�V�3��W,���h%�j����l��R8|�z/�#��GeX�-���܆}˖d7+̛э#�	�c�0�S�?�=���-��������j�Y���Su��Xf<k����N�q.�:�`�ҥ,lJ�,ՙ˷���y��;�J����Xܣi(�x4� �(��(����\�G�Sb�N�*m�g]�s���lօOt�l����8����Q�}�ó<�����B��s��aΎ4L�M$��� y��ϓm���;diٙ՜�9�|u�/���v_�8 3:be���O�2oen�\t{�E�)ҮI�{�d����ke,j�M����4L�h��Tm{}�!����L�,�KbL����D*�e^܍Z�!�eM��mhxbB�Dv
Z���K���̋<"/]��ܿ���!��Tj��+WS���r�-�K^����,P<g	����!�@�b=:�0'�?�]`�H��]���6���޿L���@��n���C~����Ѕ�1�db�N�x���:���vK<ۡz�|�cJ=��,딍r�C���t_\���5�C�@C��h+1NLd���=���
6�<��	���c_Nٞf�,*w%���Q��~��׳�wfL�]��
��ў��Y ���Y/~;��wRRof2Kh�%��]�����R>�%��o�L�Z���_�oW�)�S��9G�N����S�v��3'6g!�O�H����Hy�������4|xQ�ى:��/ˑ-�A��Bi��X��ͅB�@�V�¿�zb�u��	�{��;�T����p>;���)���;��o� �>����赀�����M��!��v�	1h�P!����M`o�s8|�
A�X?�U��uQI�
$�'9�z�Ʈ�=��*�=�kEx!{��X����Cr��M��-i�Tw�B@�u��r(`���U4HH��p���m�4�gi���!���J��� N'�`�v��z���C�B�A,�C����{J2�����7��E"r�M���jU��m�:(���=�X�E�=W�t�H�z�S���\j��T"y2}��~���\�p^*��e��
'蟥4%���X˙�Ņz�P�n���G�Ȑ�%�� ��W� ��f�|e� �J����Y�R�"m�OtF���.�Q�� c8>�Nו;����,�f ����6!M���p�X� ��7#+́�o��JǱt,�����Ɵ�8S1,�5���J_y�F���+:3��.�Ib��bU�s7c��)Q%��:���\Kᆆb�&ϩ�E�JN5��'���ǝV&�f�u��V��*��5��������M� mh;	c{�O#o��A�hc-O�?�Ì����Ψ):Q8C6�p�:��u�]�DV� ����k�p
�ȋ��Ώ�n�Ƒ�ڵ�]��ؑ�60_��T_�a��\-�*��/5;��~��q�����?X�c���1˺xC�^�Ff*�}�ϝ `&�2خ�ȨG��p6�9i5qol��!�}��3�%!��nŖ���pl��C@"�&��w�:�ZՄ���x�4�-/��Uof�,ً}p���J�*_��-�"�ڳ}���L^R��m��q-�£H.��7蔉.�8�Z��ǹu��ɑ|i�U��	��K�a�)r�߮�Q_b 8���G�!�ު�`#�h:��5yK�����D�+~\�'Ue}��}����X��n�6�@���Ԭ�̿�*��t�=���q����$C�P��c��B�z�� �m�4EIA��8)~���-�G����@�_��%�󅛧 ��u� N\ o樚C�[H��J�JYX�eW�T�p�`�}�EC0�%mqQ��ۨ�F%rϫ5���+{V�sL�SP�9^�;o��������Ӥ�*�xyL��w�WS�ɒݱI\�VG�"��.LgmN���[y�>��FT���j7��> �X,h4��m�	m&�N�#~xm�/�]�#�wC7l��vȮ��o��xJ�,?��8}K���O������yIöz��Ffs��4]A�
�jl/)����R嫄V�x�?�ך�Kg�6��+����'�w�u0�����aӂ`�\(�>0�c{M�m�*�>�Џ�Ʒ��r�������Je�*�����2�[ �]�S\|Q{���>�,�<[������|r�/���n�T�Jl�w�h�+&���j�u4���c�ʰ�f9�����	[�Nl�E��?�m�쩲��]�<f�6��6��}I�ō��Gӆ��u	,��14��Ga� ~�+.ѳ78�����<͆ު�{���K�J��^��
1q8�� �Ļ�K4\��L�YM	�~��?$w.|����N�fb**�������=P�B��G�3���Vj��� ��ŚS����[6,���o(��f�6�}rm��=(��%<#mIc��F�5��d��xI����>�2:c���<�O��_j��0�Z��ve���2̎ƍ��`/��J���/��
�q9p�ѶB��R�sKȄvj~8���+����t��9�:!�2S�@�(�<�Ҁ�G&<�ܽvD��)�� ��>$�4+lt9����n%4�H:߄f(�S�QS�y�֋��b���Rs��G�ޥ�"�Fl	��O��W_Ee���X����Z���w_�8U��(�O2�6wlx�=�o��%G�\��\{XSgg�
Y[Z׈�]zB2�$Ҟ��ޞV\u1[z:��T�IK��1�d���aut�T���ր�p$O�Ȥ���A����>(��u�h�@��
�Ъ{�񮩦+��&�bd/z��a*��t�r ���
)/<����\gD��"WD%ϑ��1�+;�%��o͈à�\��ٱ>�~p���ծ��\�]���/i� �}K:�?��C�/�ִ���ݦgoҮ���1'�6�J(�tK�1��_�윂�PS��қ[��F��b���^)���?���?���	 ����>��9�ک~�/�	[.�'.T�%�@��A��Zj
��Z]�5������$�U���}+'g�%��ՎN�j2�[�^ɿ��֦�C��M-E�k��3uM:d6$;2|�Co���h�.D����qbw&.�p��_f�҅X�'�R�*h�¸&�0�+����i�^���)�ym0�Y�n�����T��I�uX&��mU�f���`շs����C<`m/)�GF�J(\�[k�HR��t�RIG��r�R�� $��i^n
gb�⼿,UZ�-25!\~�U�������A3�ӄ�`�f�~ ��6a���<���~f1�i�nM�<<If�a�_/�ȧ@��7�j�	�l�o=�A;��ԺO���ʓX}�D�Y���c��Q��e�$0�|��?M�vSW�&���8e��T����l^�^�NL��j�M{jh�رZ��A���D���j�@�=��+pq��h��i���#��Da��,��Iؘ�?7N(B&*BH�c��dY@r�oU꽐�l���X��M?�V!?�ne+4�)v���Y�ؓO�\e�� �x�����'i$�q����hFF:����)Z�)���ͫSAzv6�P��GC�P�/�Ԋ~s+M+�6�1�v����+���O�_:�Z?�ȜB��{���S�6}c���q~�f����K��?\�!���ܮ]�tz(aZ����i�ȯ]�fD��*- �,��Q�G=���1ٛc�ޝ��E(�rj8#k7��X`F���|
*�ʤ0B��i�9��.�\��9Qܷ����hĕr�Ƨ�DQ3�%��G	D�3d��'e%�LeEq�RZ��zB��sg$��<(F�m�ӟ��JSo�WcC��� �J�F�o���2C �iś9JM~���l2?$�:}[��-���I�#/*?Jv\�������ص�$��@��Ǖ=4^lN_F���:y5��b��+v�eY����"��f-����A���a��g��#��)����;a�5�*��>T���)���P�����Fcz�ʾ��#5�����	��Z����P�i]�|I�g�>������YK��cJ��%Q,v�I��b��آ ���o8�O�����PA�)��+�-5~+�b|[7Բ4w���)�n
�l����1��J��L+�/ZW�˒h�{HMﳎ���r_��W<9B�N����p~f=�Fb�����rJ�U�L*����f� l�T3��D���U��k.l�vtߊ��t����5�J�}�b�>�ӗ�j�J
�����M29�Ȳ$�' mt��)����vwL��GC���}�e�I]�ZF7�iBW��S�ׂ��B_g��Lka�gMe� �ƞ
y������?x�}{��u����[��������8A������X���B
r�v{��<���/��1i�;��!Q6>Ti�C��*���y`N���G(q{��4�4��P!#�.E%�v��<�2�{�u"e#4�㩦�I��G�H�j�m)�$gGKc���U�V�.ٛ,�����]x����?�2Э'���:	Lj�oaЈ��!�D�G{��%s�i$��G艃`Հ��81GGn��S���{~E�Kd��R�2](�oIU�:z�E�d��6B��)�e�O����:!���`)E����7umD��B* 3n��	��ʶZ!���"i��A߽2I<�B4��3A=ea௮�@�	�3d[l�x�m�:���wQv�B91�K�a�C�MJ�M��;���_׏Xsé��?�3�a_����2V7E�)/L׉n+�fD�[V�����y�u���9[�E�;��/IՈ��[^J�>	F�+�����%�[{�~2	C-j�}��wU{p�8<�2׋�6����=�T?��9%���U����zߗ�aO� g���@P}�	��R���#o��|9⒙]c}y�v�:�n�v�Z��Z!�Hg�R*y͊��h�ȣҏ����
m�����a��y�Rn#��p�H\�����r4��X��fqU<����T���eY�����B�/����g�Ef���d�)fL����c���9pO��)Q8�������_���f�&Z�9>81��2��H"��UT� z��jU���٩g<{P[)d"-P����G}~�MMP��j��f�����{k3�2�I�r�ɩ��Ӧa<�#OI�[x!~A�Y��b}n??8
�K`L��(�}�:3��"f�i������.cB���q�CC���S��FhiŬ���^{��ErS1;^.j�\pU���n;Pk�P�v#Ne�UP`��p��#s��	A�=�B.V�>n�0q�C"o�~��5)��S6+l�^�#�nV��*� �(�~�z3�W��0�]v��'��
��/%�d��:���)�C�BIT�}�R\]XwG1����4p��Ş����7{d�_���T�'嘺� ĬU��Qk%*�=��5;�C���vi������![r���_���8hUp�G?�����y�AJQY����ڃg�D�H=�Cb��S1�n/�����;����׊&(P��Ύ�l�U�I�(�Eƌ��Q�f"�`iw�J}���rs�h9ϱX�r�8�*./�F4��H��ׁ�x��m���=Ri��W[Cp�f�4d:�Z�� ��^ֿ���������qeq�T��y	��働���H/���`���D:�ۮڗ�d�4+w,�n�5�6�� �H������{�BFy�o�VKe��Lr��C�A!�0zZS�4��_r����1wT��Ctw���:L	��>�/�v<gG�ͣ6��
@��������m�X��<j�O���BLUn6�z�JnY�\�����~-o��A�;�*<.%���kil½�܂�QC�;\�m�Bpp�y}M"�W?�C�%���K��	*�8�tz��D���+n����Ԁ�:xB�V�ӯ�?��yxF�[[W��	W!�1�&dH���@h]2��yM�L6��� �.e���UA�B*rf�KeF�Q|C�镪ڨ��F�p\qU�^�����iq���:Ժ
kB�:a�Z��D6|KڽQȎO%.$V�N�ܤv�"Pь����ףּ������t �N�!�qj�|�2��۟$����_#O$�2E:�P;q���U�5�r�²-��2t�*}�,��(l�%�L��W���L��O�B6:W�w���d4g���G˭��XeX��	�����>�Yn!�q/	�1="��t.�8V7��2.* ����7�r�}c
`��2�����0o��� ^�u�Js�^:��{��;����ܖ�e��P{vu��$d��������@���i�߇�w��?���3��3M~�]�o�9?���!'��9�4U+ᾊ��o �:��UD�cJ��+=���|�1���_k�e���R�D�޲�W:cx�����9��e�Q�i�5�-O��i�1	���B�����ϼ�_se�ٖ��l�#�	⺘�ҷ
짌�ڰL���Z��^�Q�"�Q��f��1�Y�EdR�M�2P������}H���Ԥ6��68'�z�6Ǳ�U����
ŲB���l��L�Iu����&ul���o�R��[�8��.x}5�2p�S<:eY��קT�y���؀}l�x+�.Q��R���ߴS�5��&"o�Vߣ4>JR*��E��[�ȳ�qE
����O�:�H��:D�[�Z�+l�fv&M�ӝ&����/!!�Ő�T D��9u>D��I��@��	ꩌ�ӄs��4�$g!���!���Ŵk�t�������E�����)�r\۔"�W�b%�1��b�@`by�td7p[�c�d�����!����͂�ej��$.��S���������}���M�)��jq؊�(,㏂]}�Dg�5Ԯ|z�h��z�d���Ň 7�t歰;mѐ�z@~ �����Az34k��<��n3
��kh�>sT?��E}�X��0v�n\I�y�ׂVl��ă�R�0e�H�&ݖ�����2�f�]���ob�#y���F���]��I��@��*y���SO�����Q��l�w�� y�%Eb�h�����U�	���zm},�>p���s�hEG���r�7,� �	u��n��mB� X}��^Ʈ�V���{%^��|#���&�FF�k����L���wڥ�/IK�(�jE�eS�[xG8��8l�iQ�QeV~fI!+>�%����:g?F���u@����B��c��W-
K�eյ\��8�G�U��#Z�Y� qe��
X�˵�(�J��?H� A�qŬ�cu�jr��`�"��T�X{�#^:�7��iF�i����B����+|	=}{IU�|��,�5��1t��e�k��yCX`����_�`��E:t�'�?f[4���l&w��J��^ׇ18�E�\ʂ$*ݲ/�"C���3^�yG�|,��5�>ۡd��O)S���Bz	� �4���R�����~�O�8̝4W=>�u돡r���Qp0��
�w0���`��D;���= �G��X7>l�^|���7��R�jM5�`b3��X�Z<#7��fDSĔ*ri
�E��tc���[���w��(2�N�e)���I�18_/{�o��e��X���$����Sg�|WX,�u��([D�ˡPc#���1<_��������~,a�E�3�?V�g��mz�_̏k"]-8�JY[��ϟ�#��U��v
��R��b|��_��ݛ��~���Mk���7gAƝ���c������x�T� r��b�B�O�cnʑ�}z�|��{�~0#���ݭ����	�33�=w$(}u��n�OH�W>b^%,���WM N+r�c$G�,�Ճ0t������1�+W����TF�tϡ⦖������R��e�r'������<�fh�"��5h%�3 �Ŀ�U��^��0
SU;;;�j������GFV�*1w~���N�xOs�j����Q-��3���xD�^�|���������#�-v�U	�Jr�� [�.E7�E)��j�Q��%)�^��-`��x�L���ǁ}�;�����
��X���O@�;��(	���ޔ�r��v�������i���EsЋ��n2�'�F�..�^�{&V�U�\���?�Ӿ�1v}f9u<.�H���!h���!�Z^&o�eI[!p"Io�!����0F���m�*��Bb�`^��E��cn�[�,��Nb5����%�t�r#'hs�v�3Q+�6y�@4<~�*�U�:��� 35Q���%!�iE�f�r+�t�j�[��#�IQ霎1ف{������x���ɸb�&�[�,�a��8�(^�w����ATlq���ܡN%Nƀ�L�'�Í��ߊ-������ƥ�|G���4��a1�2�U��Ra�]����p|e1��-�bU+����s�[Z�R(:���b���m�;K�\�R�{qX?i��ّ���UC��F	�h��	�b���r$H��/x�޹�����>���=�����a�϶T�xs��e����j�e�����o`Њ ~�cD��Kzu��{�����Hi��,�=��؃�ÿD�ћ% ��4K�L��3�n���}N�czR����R��qh:;�1���r$�Ū����H���o�w���j�W�d�#�!��đ�xRo��*���i�+�B�M�����S��U��6!wD�;/���J��������E���q�F΋���%N����^}�����3e ���3���f������i���TA�Z����w�kV��)N6�8��j�5����9���������r�(r�/S��L��Z�LD[�nF92,�$&�'��0�9aV��
���Fg�@���[��)5�M΁N-B�B�v�& C	������(�My����]pZ��6����J��mw���gg�/��U�7tV3TPN�cqW[&.e���%{��=��f��66��ಿ�e:O�2ܬ�V�|����c�"�[��"� 9W՜V�Pիĸ3�[�	v�>��������)�@7��'�]�Vh�橯�@���m�T[߉���u���u���HK�5-qS�A���F�nf��Q�ڂW=6��z)�,r���62����=�V^�FGL���{;Lv����x{w�R�:��Mť�f�j��5���O����CckB�J��\4��Iq���˜i2����\����T�������zw��5�:��Z6?%���YM�y�Q7"�E��NsD�g7�\����Aڮ����3/�GP.bp4]큡9G��k�R)�=��܅̭�1�$��헝�c=�S������?As��	dz��9��7y��s���E/�g�m���i��u2�FI�^2� �٤�j?��Yzu����)��ՙWџ�%F��B�X��ɧ69�Â?zI&���%z�;d����#n�b���e�ނ�8��>s��?����m�r�؄����� J���OFp"$&q��7%�]�I,�tf�W�w��|Q))�{���5��K�!*��璘ڷ�#o<�\��u����Q�$�*'����3G���B���)�R��W���yj�+v3<x��V�Ϩ�o�t�?�0"�en������O��G��1��s"���!��q?��)�;�+a3c9���p��2�+�t<����-��s��p|֟�S|�LQ�u��B��ȭ�V��s��Z�F�����HNGZX�(>�s�����n������N6���I����k�FO�2�T@S��矾g/[Ӊ�)�i]ʵ�����<�xw@�v�bQ~�UȺ�M��:a�l��ܦ�f�<�~�5y���p)����$[@�y���?w����#)��*�,���m�j��S��l�߽?����2-��n|d󐹇��YA�1�s��
sZ�3X�&���]��f6o쒰/��n�Rw��~"y?^�^� `z%��|S�D�ػƞZ["��W:���2.O��֝��f���K�eeA�D1}!��}�	Z�t9��e�nI.+�H�����D���sݼH'��/V��W#�e*����Is�����Py}��t*
�oy,J�P��<L�U&�\E�p؇�O�?����u����L�j$#�թ%�g�}���4��2wA�AH�(���VI��L45K��|.�~���D�~۳�O�>,�@aˁ����\ق���ߣ4U���2�A�$3���R+W+-�0��`[�v�v�{��`d�&�ʝ��d~o����&_�#ق4Ȟx.�^�S�j��7��Q�����P�W� ��2�֭�~²��e![qF���q� >�7:p��Trz���O�Mo?$�>�^'t�N�|&��9�p�����tki��:�n�������Ǳ��ָ2��+\BB�?��P���3gk��[7ꪾ9g���e7�(���Gn�*`�C����{l�|w������y��>�Z%`ں��1�1Ja`Oj��>��>����&ژ�^>�u
����Y�i�?Eeo�J)�6�����8u]������hp�fpgQ�n�ЏX�NHh��lٔa����V���r�<�R���|��Ҋ�($x�+@��3�y��p0M��כd�3N����g-rZf�o{���޷P�љ-�'Ǘ�?������c�}��͗�Lkb�m*VȽu�Pv�
ǃ:\����6˴�q;d{�*N�@P*1$ZYz-��֌���=yA׻W����$�0�l'h�yr*�!���yg���1.��]��,��������ٷ��5�X>@,�Y��uy����O�'���p�A�g����;��{�e��7Yz ��F�w�]�_S�1��������A^<�	v�����f�S[U�=���R��Cj"�h�	�5�n�KT��l�+�TZ_V��D�?��
��� ��_�V�}�.o,�-F��n��:�q���B�Ԥ�6�u E�~S���3�����d���|K���c�G�h��&�H�s�:��J�/	*Ir>�Ѫ���K��W��f'����HUs4�Y�y��V�Y�8�#����T�u<Dqt���
$��>�!�l�k���JhV��R��'�?��T�<a3���r��9�G���LǸP�9��rzE����*��^]d-W8�C������g�0VL�=�����X����ˌ��Q!��i|�Wm��:<���w "��@�9�r�%2�qLe�%��'-��gr����Jcx��,*�tp1�.+�"M�'U���\�4����9��u�"m,K���TΚP�C":��P�tw@���
��c��*�T��%��B8Z
O���`���La��B����:Uu�1�_��:_�<)�\�_�:R����{�f��K/�D>9:m��õ�f<�^yaիHHщ���0��lw�N�#y�S��s*�Nor��B]�j�8!�}U<�-����N�&��������O$��>�P�)��y���m��f'�D,��a�c78�������z�T� υ��ڰ���V̀D����"(F�+�%�c���&����_ ����]n9� ]d��	�(��f��1K�Hv,�M7Z�6�k�R9ꅞq�kie�!�L��"ޜ�myoP#,�+wj�d���ċRe�R�_��ş�5��3�o�x~���)��ԯ4�� �hi���1"7(�:.9�2��t�G���s�yGo����.��3��@0^M�k�.S��&�G���"ӹ+�F���oV���N����]8F����d����`3[YU$��-+��ă�C#SGI\��N�*Aa��A�ǿ�ߓ~R5�ϑ���$ �Ȓ��]/ 39����_�!ph=*�Q'���|�ߑ��7��"��[_~թup{�� ����O�`��0@A���S�p�y�	�t������������0`�Q�@T��]zu\/�ȹ�	y�m��z��%!��w��x�R<�~�L\0��_���mq�ٖ��E1��۴�06���_b�la�f�q��}��li;#O�4,`���I~����V>�c4$���XǱ�yZ�}Ҙ���l7�'�˄L����b3���oD����8V���.7���=���z�"l�{�y�dC��-s����o`!�_x��*�7l��g�m��_��~�f(:��uV��2�i��|'iDa��������e�o1̳�1�o�lk��K�)k�n���9�Lx� J�dGrI���5>EJ�m���%*剩s�aēJ���a�0�Q7�ښ�,��W˫��[�^Dny��+'@L�J������v�L�Jrwj�Z���<uL���'F,�u\r�s�e���WU��}3N�-k������3y�(� �h�A����E�c�Z\vI�y�A����8�7<}���@�0t���)�a>6��hR�Ҵ���6�	�f��i��F�]Tmμdj�T�Q��_f�\+Zpa�L�#?��Q(�M/Nv�u�x�D���tѯ�&X&�	�C�yA�^wT@��m�<$Jq�����a��Fn�@c)�կJO��u�'��;����*'�#d��m} ���[����V�Ϫ!���k���M���#`�k�y��Jg �)�����g�m�F�Y�6�K�?�I6()<�8M�S�˂�jҎ|��ܞֈg�Sd�֭��y@�Z%Tm�D���ǩ������o�.��<�%o��U��5, �'j&2����5���7ݝ�2hpl�67��IL�'2��i�]6��5�.�FJ�>L��⾦;-���Sk�Y�nw�!�̈́|G��0&W�e+�1N����ы�<:
QE�ʩ*�k;�	�&��
�����wh�`�j fD�xrD�~���O u��2ε��L���˿O���4�4o6e�n��:3�Du_(�=�F�%م�ȑ��}�H̊x(��fjo���Z��);V��*�أ�i�V\��e2+�]�T��b�O+�[F꺐A��P�E�U1�dT_�����mcZ�@��	��m ������f�KD��hmQ�u���=��Z���Zg��A{Tu>��༒m���.�"+�r i���R���҆�1"�O�0JlJ��sԪ& >�iaSwXy<�?۟� zgj@����}�Lk@��ߵo9ب�~^tȆ��-���[&S ��Ҕuz �������%��|.�&��:l���2�}mخ��5�5���H�"o٤ �h�Psg8ߝ޴K�
��g���%<�%.-ʶC�|2r���Za�w�����n����v��9��7X!�!Վa^N�ER~'ZB'��(=ϖ�2r)�u�� ��i��K�m$�v/�A����W��ͤp���1|Dm����=�Z���ذ�G����M�w-�w�.���2ox��k�������8���:MaST���(��.�������˫]�C���
���n��u{��ސQ���`��wЍ�W�e���h��I?n�g��{��i�K��8�ކI��t�f�ܚ���P�4A�\]��=9}�)�?��dG}R�˞e��y�E�V�*4k�\*��{up�@�7*�=�
��{��=���DMK��|�{�3kX?";� ����0�J��DRZn�x����@M,����F����J�4�>z:~O���sVW
&����Kr9��u���C���פf�����&�������5��p}}sab�z����2���+
�Ҿ�*<C�1���U��U'��U�l�Z���i��z���
Gd���-g��R�2}!�(���05^����Px��}��+�P���(ޖ��P�#�=LTgs�4�T�k2���v�y"li����O��T�^M ΁�Mh�A��^��E?�S�OM	o�~*�\k��oL�Ex�7����*-EA���-�/�*��$�W�W$����5�������Kp ZK���(��H:QO3��g=}��i bI�=�������H �U��G��matq|��� 0E@#����m��M^��,r�?#L.�@0�h��┚��wGim��>{�S�/b��n�,� ���d�E��QS�|�8�MN_jp�J��f �:Q�����I<;1���`�n�'���)�TR��"a�>1$�9����ʿ�U&W�щ�8,�Fr���[�B8�'���a�
x�W����6�R�Y���_�sn�l��1N=�e��55�疋��ro��OB�F��J����tO�s�Ø�$�����<?I]N�4u�����d|֡�����l�{"6Z;Y���N��m@�[I:r(��đ ��Iܲm0�ȩ�
�h������x�.��A���!�(�n喫Ѱ��n��C-k$����e�-��q�ª l[`��"�I�;fA5�:a�`�����|{�^�a�������i:с��1\���$� ���3J��aa�e@)��aw/�}2����Q��X�2l�\P
��;�����Wr:�I���T!�N=�����~ ���n��k�i�&��4%3�,YhN�wP�����?�Ɇ�o�. ��̅�n��y^��#��\��/�Ӎ9q���$$�es��f�hA�����C�e��"d�m$\�* R�o�X�x��fڑ�e$�s�&��i4~�ib&2�ݦ޹\�0�<!�;g�"o��A�3�RFY�}H�<Ek�`^b<&�9>�}T��{�ZcE�k�:���U�����rc �W���@n�:ٳ�4�K�0#	{f�`L��Y��Z�W�V�q���4��U�ys/��������k��"D�'M��*�[�����st����8H�ɸ�ዛ�ὗ��3q���A�uA��@�ǒ��J�U\����jNok����dO�1���I�G���I��:/����gσ��{R!V6=���|���B��~W������㝤ɹ�' �߽	ǐm��q�E���Vy^$3�S�5#,r�<2ey�mKy�� �Y��nU�m�[��d���q����0)��G�8qCp�&lk��,��`���m��9!E���y!�S(iY@�mʽ�
6�|���_�:x�l(:�V���c�S���q����Q퐮 (�����_*�h<:�t���ؗ��	l;CG�șS�M2������	lS0�}ʚ�U��˳B~���� ��rښ��M� AeW�<W} }��)��j�L �/8�{�~h�_Q8\�W��̉W��+Ps�q
�Gm'���~3���Ӥ��H���.?n�I�M�d��:��Ȏ`�)L1䤂�F�Q�ͦ�6��՜Xb��G�aPpI�O C��m���[�8�����K�b����KD�ؔ �2/�9��Ym����~M��?d砕aٕ�H�60:�}��������[�S�})ҭ�[z[ێ��a���	�'���'�f�I��� �Y
�|x��\S%�_���k#��� 7��ea~��p����F .��CQ�I�S�6���Uy���jfv�^�h��*�l
�ᙄ����s��w��)�Z6�T3��D�,V=6TP:��^&�]�����=�s�٠�D8=�Z��@شl���.3�ߟ~N`W��_j��S��Ue;����[0��A*�J>�m��d��>����W��b�|h��#�aq[�+�P�(`���d�y�گ,�:%�-v=_�&G�yXh�[S��dت�Z	�*�B�z��֋���n��_�^����
!jy�=v2C5�S
gF8&gAvf��9��^9���K$�-$�ܓ�@/���w�U�|;�������k�G����$><'��*K�쎳��"]<���&oUFJ�J��M�pP��;�]8�a��l�ڪ�yꐰ����4-E�V�`�ӝ)O��B��j�*ns-ϗ�_���,��3k�cT���\��-�"Cͭ}3/�X�R�(Dk@���c;)7�c7%lm7B�c��"z~0���/�m"�Ú�:�i��scx�U��;*s�\,��h���+Ș�ܘ3��Wb�1�a���=8������
�6-�Q�$���HtÊ�j�ŗ��O�EP�z��!�3>Kir����-}��#ҍ���~\�=��a��3w��|���8�/nB�3��I隻�tq�l�x�-���X�L�ō[���t4ͻ& !d:�q��j�d +j\f��#G;2�*�h1�ż�Ce{h}��4��F��s�w[����e�J6�d"#�� �[F�}���QJ��:��A�?�gd�=IA�0	�AH���$^���=ee��d�l	M@�}��YK����6�	����wP��T���.�[,�O]?�a_>�U����	��I��ب'����3`�����d轷���1��Һo��e�xz���?���#�pM��&�G������k9x�Sȹ�#lJ��|�>`Z�+��D5�[�b�y�U�b_R�p�niA_ǈ��~p��w`H'�%7� �C�k�ߑY�6*Ȟ�M�3�a�e���D��V���H�ռB7n�a'MC1Z�p�\]Oa�NI>I����12C��B����Y�6\V§Xb��_{��l�M���<Ei�U�[�;',�T�!���+RϺ� ?6v8"z�rD�3ߠu��2��R�M:�O��z˷O��n����β���L/}Tf<5�L䧙���h��?�	g^S�ޮ��c��}B� 6�[l}�6�[^��(����Ҹ���q�/(*�U䮹Y�-����:k;��֪���q-��K��wIjf�T���B{O8�}U��3 �,oTͮ�k��f]��������<���c�SeUYb[nR�E=º����tۏg���c�^(^I��� l�y�գ�Y�ؓF�ƣ�dP�����$�.��G�v�g.�5u1�3]y�8�/�ͳ���h?�G���x6�+�/�\<�c�U���B&��ly�t�W'J��t���z�I�{u� �o�Æe��r�	���3^^*�DjT Wg�4b�M:���m���z9�cIw�\^�@��<�\�+��҈����#4H�����M��M����d��f��]k:�1Q	z"�?��/�l1H�ܹ�4t��r��[ߺs��B'}����øHy��͎6��W�>-�p�zD���}���N�8إT��ۇ�x��<�BՌ�W��,�9!m�/�_l�x��:�Y�=w>
��RfJK�~q/gF�Η�şfzB�0〈��y�Q�]�,��5t;DL�-��NT{bINXC/(��q�C}%a��ͥA*�>q�3�Ӳ�H�bֻU5z�3`_��0B�gN�I��'���y����~1ut��QD�2�D�e���Ħ���z�Q��W�/IQ��9`|�7��i��6߬�-"Kݬ8�����+*�f� x�+�t��Fz�G�-����9tEDǂ~�&.Ճ��(�P��N�V�z�����ހ�ciD�ߩVP
&O4�^���1�-q�@��X�'6��u�C2��U�?����A#��J�#C$�|�Dgz�U��j�}7e��"���8���'p�ԗ6�O�/fω�ZĿ� sR<��P�el��h �:�2����I�:��w���6�̖b�V#���ׂ�#�Hs07>�[~]���� 	����C҂֚�:�Mw�e�@q�)�*�㹛�����<*����7=�0N�:d+��3��P�-����؍A�f#z�7�������� /&�z>�w��eH�p�g�m�u�����UJ��)P)����;N6��p�Q3_y��g��}�Ό��љ͎H6�'��+^Q�g5VCH������'��7�s��ubO�,�/(b�}��zx���	Ԩ�7(�i�)��`�+^	|mm������T�ZŎ���C�bߋ8�V6���r�>��,�q*}.U�=�L�!F�������̬?`�\�i/�^�4k��1䴁Ŗ`�f?K�f =��㣱��J"(y��B���v�ӱ_���/� 9!8��V�R2����@/1颮���s����\I��_gX|�O��`:x[k$�"0A�ȿv����Slk�sԗ���{��U7�*�sTM���r����Mp�.E8����F
n9]��I�C����-~c.��E�7�Y0�H�ϯӡ�Bt�s�;-��<P�/��c�����N")�+�����1/� ��=�i2���K�*���{Cb��#Y��d唀!v�h��#_;����Խ�;ʋX�J���6@ڨ�qY������rM��L�u�H���0�=_%�'���v�vJ���үu�L��I���Oq�aq� � =�cЯ�K����ۛE~Ɂ4u�A�c����{�L�Zl[g�Gu�0#8[����7~�iO���d���������7�^�@�l����7)�Xy�P��M�uć�/>2�9UUpt	>��tk433���w�"�lm+��<7fO���~L!WRjk�	;Ș8z2�,�V�U8��UA�8ˊ@0����h��e��;*���W��� �%y}d#����*3ʈ��,P�q�Y�ciz ~����eJw:�?����6�O�ā��`H[q�}@�%�|ܴ%�3��+Q�CRl�� �������;P��H�}��g�CC
�EQ"�Bjhc�Q�3��еx9O��	]@N4���0�h��K:��?�V���Ʉp�����"냫�6��GIB��.S,�XBJ&�r��=;�;\l������?���?�_���w�|@�d5���G*A���^]���22��/�i�T�|��W���3�(�cD*R��������'��G�M�joL���w�C��Y1�J�/;Ç$�߃��L�څ���ÄZ	t�����? \�th��\nw5���Sk���_NVٓ��v!��7J�X�=�/�TY�r������3�ѿAؐ�GlV���g�z6��GҖD2#5��Ӥ�S*���xo#Q�GkQ�EG1ѩ���7��q�
?�'���>�6<�/5��V6f7����1
���Q�2���b�H���F�|6$�f?Cw�׶#�d/ �g��ו[yF׽ ޼����Ql;��_L��w��hR�e�~%�]�qޑ��Z����f�/����H�
R}EWu�#{��|�|��-�-����H;`�ou��	�Nn!�������N��B�_̧!�O���ǔ�j��}����M���ѩ�xUV~
�3AU�<ݚ0!E����wF�хj���簼mP����G2Z�
���(�^�6���+Sȯ��Zz�:r���K������;�],]z���f��`UR���2}%�71�2����%n[0��Q}�-���N�?���~�DP�U�(�b�?9����Vǔ-%uC���b|c��n<<�}���SG&����~�`f�	h�L#�\����Fܿ�G���OFR`1�S%���� ��Cڶ2���HLհq��0�&L 1G�TG�-�KK2OP'�~��/�y�t���q��Rue�T��;�l����Cڵ#��6�1�®g_�_ b�{����5w���HUO8�-P�%�?,8�]^I��;y*[����n���^o���@����<��oSWK��be��K�dXh�k[�H
]���cKI{LQ �V!�'�کSy���2���aS��X k�n :׿)`����w7^u�=뚵s2�Re�qFE���H+W����
,��ᩘrL�^�� �q6���3�G9���4X�����\��� @?<��W"�mW�;���&��d��m߽��Q@��4����
�ѩ�JFWg����������.L���b�ǉ�V�4'�P�.�t𷁪n�&�f�N�
���2.ә߁Ġ��/�梂�q��I_�N�������l�D2��n���oKǚ��RnݘdO�|�(A�8��������ȮX�rM���o�%� U�Z�0�>d��l#��3q�e,?�"�K5 �ݑm���=-�v߀u�:Jqٮ�oVE%~e~�-P��xue8;J����*��5�vW��\+Lo��W�I�]���k^�m.za�>I���'S�|rm�h�Ī4 ],��P:����\m�]\���bT��>f�XR�"3�T�(�-��(+s��k\(;�3�A7��p�����kqU
唉��LXK�4��������a����:y�s�1?��h�d-?O��"e�4<r��0���t]�%���]��P��"�p�[ïȋ�a],��-�ܸf�R7��NX.����?ط�
k��j�y��o7#��f"o�8�Цώߞa|����2�T����>��B,\lx���J+�c�#A����O �՟�H�U� ��]�o	��%eE���bH�L��X��IH���Y�gفh��d 7����_�����4ɧ��SIAq�Q����o���6���ȑ,������|��]=�T��B��,�H&���xWg�<�Tw�,�Id�$�B  ����{[����&�C��S[0@��͍������9R�^7D�i���ڠ�P�(