��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z���u���<�Z	�<<�W?��i8w�Ke�N���~�	��cD0I�Ƹ-ۘ��d��Ao��ϧ��k��^
j_���{�aja�r�x53IgC�G�h��T� G�g"�c!����2���I�U<�? 5p��ݩ�L=v��L�0O`��������	���Y�uU�舻�een7"� :�޷�e��/#�����[m��(7�g77�ݬu�-85����|!��]c�x#��S� `SNV�]��_�g�q�VdM�O^����jݛ�$F��e�g�E�ԉ^�N�o��إ��8)E=���	���֫���:F��X#����:���|̆�#Zs����A���l(h���<����تGf���� ����B�������+�Fډ�VC��S���º !'������x���-�$��8aBej��C�]����``���PyM���0�m�Z[wi�;��7�eE~�Vu��4	� "<����2Z'�	אs�����N&{t]��oly��Sv���F��f��Fo�)7���_uxbz�y���X݄;J���mU�B`�_�~�$L4�������(	t��P��D04�R6���NeH1�{p�Dz����U�H�Va���x�5]��9��@� =��ݜy8�w�E�WgNU�v�j��g���}4�y�ޯ��eBŗ��j��
E߅AGd��g�: �Gòv̼����]������Mm�˦��D,8/݋�kS���Nu�����j�����;�\��=k,������ha�y�)=_Mp�����'��&��N���^���UM�wӸ�Z��px�S����S!��0�n-��d��Ӟ��3nf�s�|!�$���P�0������f��xv̀�����JHZkK�����R����\�l2D.Q%˵,�q�B#�X�ף{�[d�P3�/^#�Iǳ{>�=���
!.$݇�k5$����%ǣB��3����j�.���4�Sq���Q��s��ݹ�Q���v����Z��7���Nǭq�S���ͰL|���81>�(u��=�����e�1`D]��5����%����A�Z^H ��z5��{j��}�����%��*�ڒƍ`a�D2zmEf?j[��$��4�2V��U��}0��R�������� ����-E0Ϗ�g�VP�����2�x9(�8O���G*�y���E�B��p<������C}KA��E^/�H�-k��C�8 ܖˆ��ap��R6��}��k֌�	��a�"u��T�"EBS�]�gX������+���ǲ�Y�V�{��o�&th����9�hz�#�d��YܒXŽ��j/��Y���o����Y1���s&��%����A��0�J�CZG�O�NV�g��l���6Q7�[|u����;.ڎ��#C`qh]c�]J���T�39��d��0�eq�r/�1�ے{_�֓�}�:�_��l�3�1M��)�f����l�D!?� �\�L��6��W�o�7�+I� �<��˷��i�%uIX�A�BYc��Zih���ɋ�Y�yRu�Cco��^`�E�B�bά��L���Ҕ���˯�
2B+3��+�'n�M���f�b�iH�֝ޓ6��0�U�<���S��� }�S4�VT�0���\J4���3�d���hT�/)��ވ�T-�j\��G�{p�ܞݢI�ґr|�x]N$�#ܾ-������Wx�q'v�iN̈��2����<��{�b�(H���d�R���d�����PE��9�gh}�{0"e�YY ��B�B��E6\{�i�[=�_뙷��om�@���~j���5�]��XHj =/�تS�e���N���|�	��,��Y]��RA��&�(a��y�@ȶ���Ɩ�at�f�v~�e���
s�ML��)�H���6�|[�kD9�ۥ,OE�zw]�L����o�~��ͱ��p���\�r�./�7���O*��ǥ�J�Xk�*��
��y\���"��NX�ě���sZ �&i���r���朊���, ��^�����u� �Kʂ��W����i�dRLk�c���4,�L`hx��F�����z��}��PZ�8O0���5~	���$n�B9%/�bѨg�<;1x4�������DUQu�U2�)��[�	��u�V�s��tX\SO8����d^ߣǳ�����pxc�*� �
Oq��h�[l8�����k ͹9R0����Q>��e��g��it;˅��̔�ah��mN��x�x�!�_q�~�
��sz�n&H�u"�;)��<��)�@A*W��%�<�m�xt��[��p����� �(n��K��4,��k,E�콖�� �][�c�;�R��q��c�y�R����I�;� �Ca�m��'}��	��G{af��ߘ��}v.���UڶG�BX@��Λ���� �P�'q����	[]=�hw8XC�~�ů��\"�as#��+�y��s���f"͔�������?{���:�yFe���c��Ը�+�K|8�=�H�V�l'�l6R��;����q8Gl+_���3MqG+��O��o;@9߮�~2ك{e�u�O����&��%z0�F�tP������09S��N�(k����y0�u��a�<k����*�V�������J�Y ?9y^���۩�1�1N7]�KV�\FK�5w�`#\��P����_b���?�.�sH=�S��T��Ą�y�>^ug�ۙ�;�$	�UNr��ԌV_��n��5 �(]e��#K��&df�3.�f�5�wO��|Ӽ�^זC��&ZOa_�5��ۤG��P�zM��yI����\��>3��=걩q��,n1�������G��J[>��%+�J�@D�x�h+�r�~0������C�֤;�҂B�� �N_�X�-�-� ֲ��6�ġ�����߸�=�H���� F+g��Ձ����3�u�Nn��tz7�ɡ"3�،���<��q#ه��o���f��7G&
��3�$a\ǋ*Ya���o+^��5�3���MS8J��~i#gU��}��M[�"���vSF.C�[E'ð�Ǹe�zۨ�ZQΌ״B�N�γ�~HCeSJg�	F�ķE��2�f:�.�y�"(/������?��J��>ʠw��R
�f�H�8"�W[U;�E�U�	�a��Xv�f�g�P�tR�_8�iM!\R��=-ݿ9Hxx�k�Ԯ��ɐ�6�����ͭ�q�;������@�,���.�����֡�iCM���:ag#"�޷
J�IY���y�ƕ���Rp�nѸs��\_���X�w��G�gae�ѷu(��5�!��"�tS�������݃:��t��3��N�ݘl��7;z���o_�z7�e��~�RmfBN���qt�g|���>3�Ć�M��H�JiW�#�p]��;��w�+�r5�U�o��!�>���I-U$]�K��-�8-���>�VgpT�}1�̼��'���|4�
�
o�R[�bn����68���i$����oΗ?t�p�ĭ���T5҂�t�W�N/~f� �}?5�g���r���u���<�����
���7�U���\�|��1I������7��S�Vh���8�q��J����h�U�0 u�:��(K?"	��|#�q"�VAHJ�5����i������[ל��Խ�ifX�P�J.��
'?�7j���c�Z44�_���7�&�Ao����������Yk���Q�G����KDk���:�񔔧[�}�v���,���%BU&LY&��ks�DO	G��9�V���N��Z#����j�]I��V�q���߅�XY:�BO��]���������u��<ʿf^��3T+-�<h�)��f(��5�,�|[_�'V�Ӑꆽ�\?���Ag1�5J� c3�v�t�Uq�%U|ﰹ�]e��mv�/�_��S���,��jI��Ij��8������!��t��C-	�Ѿ:�,X����f�����^T�������c�����J�*8=���Qx��������_��.��)���^mX]&��#-ط�6m��&|k}�Պ��kRsϮ1���X/A�w<��969�e|�IG�dBQX����7�"��W������5�gcv��!����j_�'BE �Ջ��ŏr�S�;�Xo��,@���m^j�<�R�èN��^B�e&bud���Aq?�,�ey{"WTܴ3�~Q4e�9�t��";�ű:��@X�g�����o[5bcx�d��`m�:����A�n���
l
��#KB!���a^��,JZ�1�* �&�t���a���)��| �z
�-��~��Ǫ	V�ߣ�I�艏�t�k�B�R7�p�RЉN{�7ͬ�*�8F�S+���jL~k�O�a�iYHK������`� c���4�1�$d�����";�P.Z��*��R[W���9W�xO���$��4����M�_�o�_t�:�(���-�$�Jיޞ+���ڒ�:8_ì�R֧��	�=�W��[� ��=E��Ԯ��ڈ��W'L�K3�	��PH)$H�9����s����E���()�vTӄ Ƚ�L�!ڇ���D׎�V�8'�7m��5��m/8R��(�`�"!w-��REn�ƙb)(�ъ5䘟&>�s�T�l�������Wܡ�]��tf��Q�	����>}��i4{S�=� U���wٍr��\0��<f0����[R��Y���+^=�d�=Ch��;T9�o�I�I���F9��m�48��W[��;e�W��D�ŋ��̊8h��h��fQ]#v��C��<�F�^}���c3'�[�g�77�����M���W1��
����-}��ve��.���Y�� s����ͫL�\{��s�\��;�$�ӡ5����'�圠�ד��x|�z��WCC�S��2�%�Il{����
�Q�\f�C�"8
붑|^���k2Χ�.p�lDa �X�H��h@#���Μ�3VP-����7:�*ѷ��E1�	��l_!Fc�gB��c�@g2e�vd�ݸId���FX(������L��:�*	���^�@�,V'����� UI�~�I1�@�l�-K����d%&P�2�w�|�C���R(c�\?�@| `Y�e�x��q���쫲0k-1�Q@KB�"�l&�Gy|��%W2ehٱgG�e�J��0�D��R�4�^�s�j�F[�f((��̟o��/�X�c��	�u���1'5�"\�2(�T��([_1���@;O/�"� �c�+1P��µQ�H������Q���^�=�?�u�F*io���5�c����\L[�h[�X9��({���U�P_?��T?���@J� y� ���`G�}/�)X\���`!s/�
g��l�5�^Mj����ߛ:���C�~�T��$D����k�jYv�v*~������i�=��,�-�����	��2�auTU�S^w�H�
�[��.Eq@y_-TF��ri"�_��ɦ��R��x�$�K�ij���?~r�������t+{��ѿ9*��[2� �_���!'��FrR�̜��T���{ME��b�d3yc@!7�ϕe�~Ǿ"K8Ǒ0[^SX�O]�#g�Eʎ��8�cMQ�μ���V������U@MKW�B��j=�P�~/�������m����\�2h�GiB	N�����|���2����rJ�nL+�;���1��Me
�&IɈ*�G�}���t0a�l~E��,k��O
�ĉ�,�\���ߢ=|�9U��ى�|����ؾ5�)
4�4��:�/����;@�A��d�J˼L�懡d���f,�*�OJ^�;UTC.��\��H��H(��(��'�m�ADt����ߓj�JǗR쿊F>�޿����S<?�.�ª����Lh$�L�`�;p�b�I>��ߛ�3��Ȫ�:S(J]" ����k�6����Rh��bk�)X'�g�	�ѡn����ɵ{��j�yɧ��%a}۸����|��u���t���1�x׉~M`�T�P����ԥ�L>L�W��¶d�C�C$B�����V�:�~�W>[o�$�k�zE��ʈ%&�dĽ���=�sNLl�4lt~7 �w&0u�$�7���XiHG�TG!BV�+*o��)KH1*`��s�����m���@�<ba[��	���a@�b�چ�c��׍!��h��}�Q.��b���ѿ��QdWqvr �+x�T�W{U+��f5Q@�uX1�u�L��U%�gq�h.�y־���D�u��y�~����}��
�-UB�6GϦ,�<S7!%x� �5w;�92���Q��"�9p� ��f�s�!�b�

�m�舢���!p*G���uw�Z�@�dU)ʎ��'�q�5�J����=�+uZw5���a�l�&�=c�v�Ύ3B��?"A�J6A�z�E�Ja�K�^EL�IsS������kV{4���4��@�]�͗,�6.,�A����JY
����Kx��WJ��m�\�aV�G*ZLE�+���af���+GP��8�Z��yNc%a�)��E��5iVTI�����A���ו9���#��5P+R42}�]@�#j��Rk����	�����&6	[�5�q�A����8k�d�}��`������.i���s�X���z�*)��C�X�{]�2��9.�&������0�Sp(:+���Z~8S��E`�sV��;ܤ��S���]��q���Q@�`jorb���݋�-�#�҉Ч&��CpR���k�azґT�݅j�r�Y�2��B1����}�?:F9�8���:�>��&L�r�s��}�[��U�g6�?"�h��+�d��#������=��
-�m���>�<��&�2�G3򵯑E�b�xl-�j!Ԛ��_�E��mnh�� �-Y3S#����ZBَŽ�`񷉪�2�����/���Q�?������x��ޡC��4�vtw� vU��tQ����v,V@���*ƺ���t ���	=/� �g6E�>��Ç�k�n�����gܛ�c}���?����Q�nSZ���p|dᡊ.���e8�����xW�����([ ��A��.hO46D��/ꎑ�D��jN�~�;��MWkϫ�S��:F�ە�P���Z��3�<z��Y�1�_��{|�d�|*����LË�8�?��t�����Zr}.��_��;Uf�`+�c�;��~\l�����X�h���`�#���c� ���=g~��R�B6�?d�y�m3�xx1�x��6���(NK���=�+�@PP�xM�i�E�ځ�i,)������d��RjUzB��t�!�"�h����56=Pϡt�,�} �g.���x�AX<��

�|�RJ�I���� �\8@I֩@m����Lh�DiW��0;=im���y	NǮ��/j;���;_[�.|l}J��u5�,�GuM�ˎDt�"r����uk�,����pl{L$�J������6�O��{J�w��Alj]	GY`{i<�`���)>\�2��XN��ˊc��D��6�V��\j���&����5�ް�����+ABUS|Z������n��#=���K8j|#s���T}̘ۙ[(���F%��?�)���"YI����w��֥̒�`j?2t,���Zu��K[&����H�tÝ�~~)�y��\�R�W\4]��h`rBu�y<����A���v=ȘD܇r]���遅��#�#i��VV�4҄]c������v�"������=:�3�8��3�|����1�>"�`o,(>�7A$=ū��bt�t��`�Ov>�\t-�8�b�������V߳s9�w۞�y��Ps)�m����s��v�����~-ɡ���x2c��x+����ͻ�<9Hw.���c1�$�Z��8��{i�*J�6��T����+����N��E���\�cS'���p�U|O@X����C72�\ŋ��F��ϊ#Վ��CinzS��J[���<��wnf��>3�p����([�"X��}���m���Z��I0w@c����A|z$���J�K��k��R��2���T)�܂���5��](�
��*�࣢ �ߟ��d�E6b�d�����y��6$��Q_-���)����F�D�G�rI�m�_�'���\1V?���DЩ��ǽ�s�}���o�m��j9�2�9!a�@��f=�(�Ps� {�`�:���&I�yʤ'e7�@��|Y[�K���	��N�a�E
t���ZP����O,����ѽ
��m`����+y���ś.>w�
�KP��UEm�Ɉ#��q�;�д�E�gu�)�����f�j<}KM����Q�fF$Dz���s��3S��[~�t*r��E�xMv�|Adr�x�w6���ݛ��2���d��%���
��`Tjٻl<��FH�a��y`�Tz�Hf��@q�T�����tv"U���Me�/��.p�ѯ���#]�Ԡi���§�дCh�6x�C9k�������k`Ħ�W��jp��2�% ��ժ�uW+,g��G�r@���8�y�`)��<P�-w�ܣ�Q��g��3(�x^}��R�&�������o ����jץ�T?�.	����*����~-2�6r
9��#�XY�O��C�'3g����zuq4���(�/�'L�"��|�[�G����q�S��*�%�� ��o!/鹟�	s��r�
���43so�+ٮ'?a��T������(��u�'|�|�I��A��r��O:p��7X8/���l�a��g�#.9�~}<3)<� �p��i���>3"G��Y��@�I�W������'gL�Y��T��r�H��x���[�R*��/�G��Q&��g&t@������0H���ќPlH�܊ ���")χI���죖��'��U�)1ѿ���z�N�~���}��K�{�	������m"��3ގ�bΪ�@�HrI8w<�KU�̱�����c���h��(�5�IG%�(�_͠��xJ&�����I>�;+�߯H�K*�Jrprs�I��[&�u�ƪ��r��}���X����:�ĺ��)}3��f/TF�c��O���ܬ�ӂC��Vg�HK����c\<��ٸ�U��;w*�L��Z_�C�Iϝ�%'�S���k���20@���W<r�i��҄��a���Zt̲ԃc��s�1&?-�!SpJ��rg|��$;p2W��jַ��5P��{�������'�x��6���ֹ�<�;ON�6Y�+Yy8���j�U����pD���˭n��U*Ţ�'����\sm���3h+F�횧~�Bk�LS�3d �<��
S�M�D��R��|����.��<٬(����0�!��Tb�p�`پj�b{�"X�D�N�\�h*����+��)+�P�-����`�"��4	�z��t�I=a"�|�~tv-@�;� _i�j��#�m��_����f_t�	��&�ůH	�-f��2 q�Ɩ�l&�V��-�����v��U.�ezYn,-�#�R4oȎ:���	[�/�O!��n�1�
���H��qyh{����@Ro�NN(!E��%�4S����$�a��>0y�y����i2��t�5�PI� ��5��=�V=MW�gP�r}D���,4E����
5N;Q8���S�N�J�]�����~7���3�/P�x�p��HX�A��DP�X^/E�(�����HLl��;1���xܸ�/'����D i����?�6��"JD�A�?z�k�C~��AG�U�]#�-��|��
�K��ʎ��B1+e�e|Yӎ�m�3���t��=ٌ�d1��e�[{Mh2�N��y��N�>�'��$OۖӎK���|/6��G�Z�W&cJ�E�>��`�� S�ZF�����;���FL�dXҙ֩��1!##
�c��d�}�9GȄ5�'��1-��w��	#%9�io8|�� b��-g��KQ
|?K�B��)"��[���&�&䵒:4E"N|�8�����&_��_�9��#�vt���dZ74*y��A�	�����rEI��/��;l�.4Iˮ��`���s:�\m:V`�/ءI�����%t�&��dc��Ww�j���U����Y�	n�RΎ�ތ���sׂ��ĸ������RC`�a�]v4�����5���O~Ku �z��j�FZ�NSh;p�i&�<��޷�Β?���x�YF8��M>CJ~y"�b�/��"�;�S��
�Rq�ɨ|�t���,����q)�ز�|_u��7�zi��'���%7���t�5��=���^ /���pG�U-�y+��^�5�t+��AP���( G\~t�ܺ9:�Cn�qS�M/#���An~^%����T�CfG
�j��[��Z���!�EK]�O�P�ɠk�����f|��V���JSjء���?����겚�����/`��Qta2�d�.8!��3�YR;`���bR�`��
��p�r��0�z*�6VW��������������,J��a#o�G'$b쾲��h�<��wkm&��s�j�|Y�^�_Ejv����]%���d���&Tڶ�v�P�JK��`&9�#�,ԑ	�9,#���L�KiN&=�\j�?t��`3l��K�Q:�mA���_0�1%.ŗ�f4��K��ɔ�(�*�y�dJ�P�d�ƅe`o���m�J$`-t|�ڣ�(���͗���v@�i�Q��c��ExH[
�`�8{U�6K׸���Xʬ�~$��z�(af48\'�6��T��lT��؄O.cR�42η�+BČG�E�'� N���]o�߸>�5\�Rf�@z�����GuW�:�1�!Ww>�;�^#���lx�Qp�[+P�g���u:������vB�7���LÛ�_�G��f�6g����)@q��$�����Y�.p����������	��׹��y��݄MK�mY[mp�X�n�L����KFP���L�z�ғ���A
�|h0."���J��Ѭ]���]K��.8U}�	��W����!�^2Eٴ���ߖP�,A��h���v-��+&;J�mf���5���0O�&w]���*�=�p��G�d�7�����{sM��m�w�e,=[��	M�(��ђFw!��-gL�F��T{핔��u�`z% Ub�Ҩ�xT.<�*�53�Ls��P�Y˫k�Z�4�����8�ف/�Q�U�G#ޢ�<�Ss.���"�a~b�F�nqɜ��$�^n�gf�9#������A��hJkA�c�[M���h<G�宕�U���̐�psOP&l�`��U s׮��`̞�LD�LW�>"0º浱��b��o�&��E��U�P�����[!A���Ng��nL���E��<|��n��~T��� �wT����}~�oHH�[	��Gy�č-*����rG4ŀ�7F�h37�6M,�����u�L~׀�JIs����>��n���Â�z�d�����Ք.�>U��I
4����q�p���"P7a�����C(Z�2(�?$���PN���)b����2p8w�#@/A�]eL�^dW�E�+R�Dat�gִwk�5�ƿ�)�MzPNRo�"@���R�H ۛ�E ё�<�)������'n=֣
h��K��鰒����]:�L��?�Z����p4�Hl\�g������/��	�I����*:�N뿇��H�RKȍkDv����%o�8��b��Tі���p8���a11#@zME�"C�{�9ԅ�M\X�
�fus�y�lKz�!����u��gՍ�?-���cI�H�_ܛoè1�_��&ܻK�l����d�?(�#K�,�K_v����_�"���:���w��9� ��*�$��4z�mqh��i-��?��M��J��7{��pN.&���� U`C55��:�k�w7�Wz�(�q�H�w|6$�sa ����8#eCjt�xOW���N�AAT�71.C����C���ch���X��||êU��aM}��3hn�gס�1�����F�I%���U���C)25h_�����m�`v�W�]o~�$�ݔ0� ���+/tE�"���B�a��6�ӌWq���Q	F�o��Ǯih�aBݝ9�� ��j&ry_���A�-W4�36C�������Q/�J*���J<�B��m���(�����������۬t�v�� ��x���\(��é���2E�Y�$:PՊ?拿�[e<�T��ijo1GNGm|�k���]|�����B*�C�ç=��,@�܍�[�n�ϬE�1}����}�P� ��D�Zv6a���]A�)o��(P<����\-�#��-���P��@�n�I�.�����R��L�y��(r�Zt_��Ł�+Jt��Вt�z���Ch�Bb���b��i��Es�F Ks*G��!�/Z��?O:4g�����a9ޯY�qq�=~R�-�Q�X�mqT��w�[�}���Et�ȡB�����PǺFv..R����?m6��Dl�D<T��gU�
,#_ˀ3�P��K�dP$}v�T���m�s����v�c�e�D*g���υj�]:P5�Ў!�Ä	k]�:_ �X�����BB��7��᫂#�7���{�z�`e��C�&U��ʰ�xTȧ�T��j�)�B� ����A'8=���6�b�]�I*�A�NzQ���u�r�$����������"�۸~o��eT�d���~�cA����2�/��\���:�{[@���<XG��P>�Re	�SJ�B*���&ԯ: h���~~"ь)��Y�h(�B�����V$���Dy6u��'	�s��d/:ٺB�y@�
l��-7�r���V��d��������]�uTq�a�xM����g������^� dl�n�SӯV���./�a�b����f�Bm�u9�����/��2�;OqsXchO�I�#[�^ʮ�X��������K �����gO~C
Yn�L
�,3�+zp�%ZM����L��k����L���W]�,$q0,�fj9��0KN��k[Ċ4/EI3g|:�����G^L�?�rA�ʻ\�3u]KP/��b�Y��:o��=�>m��,?(N�MP�SC:�
�<�j�-�_!Y���.{������KȪ��ҼZ�E\8["O���f@���
���9��M<Y�3}�6!�����D,���]<�C���o�%لV�_�1_�8b{3i�,�$.>���ݫz�[7ga9[[���X���(����ف�Ina}MR��d��I-~D�1��	�N9�gX���5=�!��	�=%h����Ѹg3C�x;1�0)E��h?j�R1��ɟ�
T��Z���al�Z��7̍��x�H�ݖ0H(��w ��'r:j��nǷ�����p� �ƕ1�c�s'U%� ���L3����r�ds�����;�'Ik�O�K..C|��Zsvrws'R�q�;����L1b/�\d_K#���W��r�+m>-�z��$Wԫ�co`�`�*�R���d���NJ�h�\�Z��m��ִ�[b�e4��A`,>ih�k�+�׃Z�էZ�<Z�W�ˉ������J����M]�/SSsg�1��?�*�d��";���u��������#hE�z��!����V�o�����L �-�`=^�Cf��mO��b=	���C!�������u�5���3szL�p��T��5��E�K��HJ{Oţ`DB���;Za���-�]?���qB�G`&u��]K�9���B��,���T���g4���^���Q��6����g��	���U7�� iT��֊�FF?$:�{\�������\]���tb���`��ج��#�:P���6�3�b����E���J�H��|S�Hy�=0��ӳ
k�O#06��@�$h��oe ݠ��/T�ț(8 �Рm���B�N�V��^'@���/��5xD�qx�~+����
X��^j=��q��ޚ8�be�h�r�r��V���٘}*�-PԠ���z���j�GK'Č��s������ʡ��a�_�	Ę���㙖O�z�LM����K��L�Z��Z�;6�zB_4-ݴ������|��_�T���Pk�̎�{��l�uf��]���+�wq6��b�R�C
��j�Q�n�V}�����}��iIT꟢2'p��u�{���wb�B^�{K���yB���j��h�`+�0SѢ�׾{qI�t4w���H�I��[m9L� ��7�T����}����J,��˝�a<�-:�iF�3�'�
6@׼AFZy�1q���Y��r=1O�3(Q��@A��୻j�����G�2�:��v�q�
��P��={�7�4)��Ö-�0��Y(�)-o��O#��qcQ�@��x���Z�F2[w�� yFźj����#ՄE�����v��Wv|x�m'��y-�#f��0�.�Y(М`���b1��V���O�q#�ǭ�U�����3�p��"P<)��2vd$(��Љ�(a��|K�L^�� �e!fݏ�t�N$��~
K�`U:<'*?���K���e:~)N��m��f 38l�����Ͷ� S��՚��+;9s j�6����+�� V����WV�)Dmj�J�Ug ����k@�Q~�����q�kՖ���d#�W_n��}�-ČRZ�?������@.̘�Ľ�"�z?\���6�-ã�Y(ջ�e��M�5̰�h�'j	��A��AjoK�N������U�|t)̷e���n�7�Wś�d�D��d��i���h�c������B�i4��t�ߡ�	�5Q���9�,1�ؒP��ߕT��˄k��� ��_ݥ��䢺\�:�kI��ȴ9oh\�d�q��#x�.�.:�t��,�0��m�m��6fQ[�Zd�z����U˲�W�O#�h�и�V�o�ė�yޜ���n �ī|0c-a�aO�]�\�y�O��n�A�O�>��H�Cy��w+��(^���|����eA�d�ʺ� �����`���b}V�7]��SZ��Q<^��3?��v04KSǄ���ۇ������f"<;�z'�O��b�Q�0Cm ;�|g�4��H�@�D˥1q�R�t�%�4{]O�C�����C���ʿ���\6G��9x���P[�pe-qJ��J]�R�Y�$f�Xr6� 
�0%���z<Lj.�ɭF҉Xg 1�`#�M��%x�Iq���t ��}��@}wY�ҬG[��n���7��}t~���P���|�L�\��tU����y��X�0�&��z
zn���r1��lW7�1�a��*��]�f=]����Xw�#s��_G��$J˧�;�Eӱ�[�-�]ڜMbr��v9Lh"�S�o��KCR5���L�R�:��Ob(�٪�R���)��w�C\��1SƸh��^�Qv�U�O�}/<����8�I���gZD��}��ɍ� B����>tV& �$Qy!���P�0φ\SN��:z₡dz-v����bȯ'�a�Ba*hq+���.����GTB��ñ|i���&��C+�>i�nʾ@m���\2�	�6%E	"���8/О��C��5g��үL�e͒ ���-�D��^�.��������d��t�!���8����xr�v�k�.�v�p�<�B�?aބ�iCωL���p��$x��D��F�5�ጵXȲ~�'��.�0L�C(e���}�f�����������\Ȱ��Yy�	�ͱ�:�n��wu&_gQ9��N��9ihY������>�o]H_�z��W�9����x�^�[�u��:6�	-�
u4�f�� &oux�#����YX9v����W:��"�����m޷�����[�낁�<�F��XGL���4GY�|��dI3���$ �:{N9����P}��{z�ϓ�� 8�����lA��;C,��D/�Y�m{�gW�nt���v�^G��v�W�/����	y|�]{Z�Hѓ,l��}=Q�V�08×%HS�$��'�fk��%���D�'nCŒ�͎�X�c�,�":ے�5�T�䠀�nB�1.93e�7�v�bM4���8{43 Οn(���K,\_�vp��]�I9���[&_������B�$:y��>���񏍉!{6Y��ĿG�t��׌g�Z��_���rU��/
�
��z�Q�s�S��\}\�V18�����EQ�|ZE������Dy��;��p�ma?� �M`��U�R�z9�l�X=�P�xb�U�������_gk8@;�jwL�w����~���kG[���وsɷ�WT�8�����p�"3���2f�F�%��t7.���ƅKU��1F�����#ZL�Ϸ�"��o�l���x  �����5�6�Ւ_�uT�,"Yv�W"�!H��veH�����y���gx{����z�[�V�(�"Y�dز{(���_��s��Z�0��ޓ�<�s7�+��O� �sZc4-I�H$΁�4ο!P�Pq���{��3?���ȂV;��4/ah]k�L#PFz�8�5��/�u���,����,�c�$���Α�����1�:�1׺��(;F���{)��oab�h_*Whhɢu%����%`X�%��-��K�� �:V��06�]U�XD��N��I��'��p��a��ң��AK?0���ë��%�d��=��O
���p�7�;t �.l&A�=�E.�&:UG7��l��<P5qA�A��7�ܘ4�{K��d;�'A7�K���
��;��0?���g�61�E�)'���{Aс*L�@���`�ԝ=A�Yg���tk�NP��%/D��tpԚ��[	�:X���Fϼ�)���=I��@������z�ؒ=Dj[��؟�NC������R�����=:
��|f��$��(z?7?8e�&>E�^�5�ם6��+����š@���������E:e������������f�����Cu�?��U����=X��;K��� �/_o��;EP�D��hB��¶�[�gT�e��3����	]MlֈT4�c��m^���B�U�_X;���]�PT2��j9~z�:������h�Z'� !(N(r�zT�w�0p�ܺ��p�~9�;���)����O�ͦqj���IRH8���g�\.]IcE�5y��.��_�%��M�|u%%��k��;OJ�6�u���x"�==f�K����o�k������^�5�.�\���m��.Cx[⡈X2����=R�p�o�䣠⠙�����p��� �MC���J��������͑��J��.�z������ҋ(�>�s=�����ȝ7���!�Gص�\K,Eo �FP�8��+�w��&Ү�z��s����٦S�3'��"'����0ri�N:���(���f�j�`/x*C�ˣ��y��p8YWk����MSy��R��5�V�U,Ěiȓz��a�pV���p�V�NU��v�Ը�t�	T���c�����Dw����,�{=V X��"�0�D��_%���M]�'�^Ջ��!��Ld�U�	��|4-�eJKOE��$y��R���� �Ԇ�#b�n����]^�c���d3�Uo����zeژi�:�qOL�L�q�ˉZ��l��&M���&�jf���u�aЊ�?��� �fP�.�:Vd�9�z\p�Ѝ�y�y@��)T·�f�6I��wuE	m"�/�񝎞���C2��G�:@�-'!��Z�Wn(�!qa�4)un٠�֞;�܅~��k���e�4��,̚䀠@���y,]�*m��h�B��ҟ@n�o���>�܃c�r�k�����Q����Y�~�[�*ɭ9E­i��G�Y��Vu����{��ob�x�g�$��_���a��T�Q�������ꚇ#͖|��?�,��4׾8ڔbU(<:�lOU��w�#��
�k Jݓ(���U�ZM��a>��3yF@�����n*^c����(i6�4Fcsf���v�'X)�������QPҒ�)��u:Ű���jZ��!��>L�r�,�����֛�i�'����S�u�yC"p����Κ�ܝ��^M�-Uk�D>�N��fe���`�Jx-�"��B��0��W,� ��x���z��-����~�0��Ю�}<$������W9�>�#��;���PN��?ssuF?��*����m��(���&C����T3+=k����[�����U�:�(J'��� ��4,�)���\*`TOY9�lW����`��9����ú�O�^�|D�����t[v3E�C�S{ad���M�D&�
�8���<§"��^�?�PF2��q` C?�:���d��U�m4k�O�R��,%1=��qڿ�!>��Y�M�a��?�2��<hn�@��ɸ��m�L^r'�ǒ�tcC�O7�/��J��+Em8f�=�4���J���n�t�L�2Z�i�Q0fJ0R��.�`1���5��oa���	Wlz�����G(��@���P���<��6K�|)�C��w/g��3�g�svZý�jr�E���A
f�����m���?
�X�����p�Qg);���rA;7&J���KY�!3,�� O"���Y�`D}8�_���z�#	ӛ���nl��"�Fw�y���:��Y��g�{�y���!N���n�#W�}=Z���Q�	����se�H�h�e*�}3d>]�yU�����H���Rc9�e�XD^���t�[pⲢ�q�3�c_�hx��'��Zou�`��2����hI��2�W-��m/�WyO���$\�&���,�AG�|x<ϋ	��L�� i
Y�ř(�8��K�~�-���4j��)�t��[���5����N'S��f��>返�l�
X�̘��³��'#�΄�C�r�k�����E�q�v�����5h�����v��c `4�&.����0E_�d��2Z>z7
{�����G��o=Z���)Of��]��:�<�Fq��s������6�;�9�~�>s�}�����b_c{=J���T㉔�<k֙�Z=W
�l��6�ո��TF�|���;�c�X�LW__,���2�|�C��G�8x���k�J��v�<����[L���@ ���m$���ǰ 0�6:�c��Ŋ�-k}��z�/6��u��_&P��6��0�ܗ��a�$ &W�'�t*��&����I��.��(�|U��oxڹ�Ʒ,?fn�&�06�P��Dp��(��n�J��A�t,�}�X���q�\�ـoI�a�s{�}i��l.sA��ܔص�M������_�=�[�J�(�_KM�\�'�ſ���Oib��=�8���&�*H+n=���~DKc1KcI_�BQ9��a�ϵ}U<�ЧJ��_�}��&��ˀ��s(����#5`��l�(9�^ѴB���yrÁ�=`R\�!��)�Y8��ݔ��c"x� �����/&�x�F���k����;'j\5:�9���	�V��`|�s� �dJg39$7bd�1��0�@I�V8����f�J@����7�7�(@K��	�d�����SE?�H���c�y)V,)��'��%��;�	@r�Ak��6����(��OB��z^�+7�&Vy� c��	ҋ&����d��1���b(��2��\hDPKq�^�]J�w�t���g�!c��7�Cg?�e[B��3l�F��
�T�FH`ntt&NݩWU�_���B��3�@}n�V���eC4���U�܉���	z*X��"�O��3���'`?4�HGU�i�g��,�����k��=�u���(��<���� �̀���8Y��ZX��<���=\d��G�a\<��n�"�T���b;���\���{ZX���Ӗ��ڲw�_q�moǤ�|D��1x7S���a��@
�[�qo�V]����?��&� �$�qo�C+�]y���pC����14�\Y��{Z^;DI�kg�K4��!C��XWU��̬��#�B#�'�z�x�*����+��t�z.F)Y�d���\ozY�D(mF 6"΄\6G�I�^��0O`(�>����$�X��
m���f��X�:צ�C"��:�j�nzyt@��@��p-�����)z� ϯ�Ŭ���Kp���|�CQg4|b�(Gᦐr�)�����F����߽��ꇢ߶�-ۀ�r~�U�p0��W�<�T���-'6�{d���ū��V��%�FtX�{�LO�j'uZi�x0�^j�5fn#��2�P��0kI$4llԡ� ����N�Q�A�&��Uۮ=r���HF᳹�8��:�Qb�Ӕ��V���䔥���R��p��\|�]�H��ЍQe����z�8�5��jF/�*'B��+�H<���+a��+����1�l�p�q�H���{5Z��PB���9�&��z[-@��jɱ
���G��p	� ?eo�J���N=gG�T�ˋ�׋�����p��0&w��G��ȲJ�)*Jh�?�9"���_ ���J�B�R�Ԥ~�=�D�{��f�� �he;�F ��@Kml�;x��l	�-����R'���� T& ��oQ��uk�z�B���F[5��9>M������s�^�Ы��̰h�d�?�\Ϝ]ي&���̦ά�O�1��6^��KS�}��C��|l��N2���39>x$�3ސ�y2'Y)���[��)�`r|2P~�D���>7��,�۩#�g�Љ���Z��O�۟��Y���ۣ��J�EGz�����j�����}�	���"�����$V�0r3��)Dq�ȱ&�2�N.�F�|�YT��e��NbP?j3O'�o�DC֥+��Qq)�Bo�ɉ`W�j���l�;8s��)�x)0���|��)�lD�ʃ��� %�1��I�u���0	M���	��ͣ��(�XN]�&�%pl#<��h�BMNԈhJcR)�ҋ�rZ[H4�o]�dc�t$��7�@-ߖ_=�b�q�
@Ҧ�h���������o��T�}�UNR��%Z5�HQ��A�)�zY&���+���eS
>�X�ǌ��CI��L#�Q��3��5���rz��;�!���u܌�Hj(�[�zJ�*bA��}��(�yba>C��v��[y�xw�O�`)h�����>Ak� E�b�y�u�[M�G5�(A�2�����e�bzkX�/���H#��k�*d[B�T&x��}�L��XUa��9ٙ��������M<V�?�q�lZL�����E����!MG�E��.;��Am�_��!����_,,*#?>l.��k��:�2QG,Ü��'��M\E�o%<`��H�Ōn[r��yf�#ץ�9�R��@�g�g�ly�&J;�,!M����Z�������r�T�[~��.p�4Ƅ��'�0N<-��F6��\)o���镩��2X;�B���<�PY^�D�gQ-1~�DX#"~l�('��_u'U'���]��KV�F��H��y���8I:2�`#I�k�G���$���"��L8�/�(KVfi��e�����Fwd�0�s�yШ{�;<-4>�T�vf;��E�3A�J���r9�J)�ZvՆ����	QK��1��5>�$c��i']6��\��;27�Vg1�b���l��E�2%U=�����:�SF;+���{������f��U�:j�i�`p�L&$2}�jwG�fH�������&e6��5�R�����,kG�,��*/�� ���&F�-(Ty͜&�����ERm��ĠkO9O�Ϳ�`xƍ?��h��.Y��Br�3�=i��O��Fi�S����H���F��q{�,lX���A]�y\U��"���W}��R��+�������,�Bm�y�T�y�%��56i��Ke5�!�7m?��B���W��M�em���W>������|��3�(��C�/���akV�%�=�x歈'�R�*Bvͩ���+����,DP�0�9��b�.��K��*�j�kllt�����'��k����A�]8����������o�S e���s���3�vO2��&��$.��Ej������v���99m�+6���Z���v�����3�;�A3�V�0�h+5�j9d��2���c��.�p.5�0 �@�5[��q8Eo]�ߩ����"<t����i����ii�H/
-�]j�b?��ab�z�W�n�Yg������2���_�0��B��kPX��Bӯ��-�������i��c�B��FzoV+n�
PwU�~3 v�u�F �S�1q�Q��W���I���������W���w����ᒂ��s�+�s~�gHk��C+�.��"ac���ݑ_�nB��#�+�����!ZP�٩]ߢyijx�J��N�<�z�?*oL"��E��_m���Q� �B��7�m4��������v��b�L&*����Y"�v cm?C�O��3^TL��LX�.�Wa�� ���É)U][��f<��s9���v˘�淎�<�!�x�D@��`Wk�m+��b٢h�A6�kd#m�l,�$dEc��
A`�#���R�X<�G �F��iC�ܸ�|��_1�����ev+� �M�1*6�;�.n�΂j�b�V>1!�2d2�8j�~0A��6� u�7�B�C3�^�2xƤtδ��k�^�%}��ڐ����M�[b��h��D�k�gt]mښp]�SV�9��
��`ǉ��V00�X���E��vU����~�)9��/6�C�e�"G�#���Q��;�����h%���?��T�oƇ|Y�,	f�ٴ*��=6�~���emr�R!�N�c�
8:k����
���E��7}�_*�BRs�=�2��c��C�|�f��\��t�����~��f]&f���_dM�E�k:��W�7e�8&R`�V��D:&�nE���g���m��#�v{ڗ+��,�z},�8zS(�Fp,0��4��D�E���1�nc�ԭ�~���}�~�h�Kța�9�f�r٢nJ_H��~�V����I#?�7�-�qM7m�]����Lz_nbt��t�ҿ�<��E�	o��Q���ߓZSǮ�I���z�O���2�{>��A{�"��\�Ԃy����<!͕ƪ�����fő�EzG��L�]��;��(�5�P'���Y؉Y�����|�A�j*h�P�^xͩ�x���gR��Z`���x->���%��I��-H!��w-9���jr��>K��H*#�='�E��r��9~�|!F.ه����k����'J8`U���sl�Ԍ����cc�{ѣc.��YJ?u��{�6������h����F.��ʥ�/y��K�&�x����'�2�쫍��e�褞�$�]�۵���;Ft��n���:�����q)�jP#s�&�u��H�8p
��D��M�?���9J�V	7���&(�,<n� &�0�xή�w��GCzkg��Y.�"�E��YW�X���v:��2NF�̎��P����	���u��:i�qC8}��~Y�ORn����9R�o�_�,K�m�R��Q�8�(���:�[L� �=���+!������	7J�;=�Oȹ��V4L]��b�����-�x0`l�7
�GZ��>��RԸ%ωg�a�0] y������g�ϼ�^@/%P����Ƨ.YԖѯ��q� >�c�~E�Ц1�l�O��2$��I>�3{P����u?�J��z���i��6=��^�nf-
�hfy�X��=��C&��C��9�Z��vC����E��%��������e��e�V�#�M�G�t��t�CG�a
9]	�-���E�XbA�jB��P�f��g�"_�B���݈hU�!;e;��_��Gܫ�XՋ݊�Җ�~ƀ�8��®�V�6T�'����`��>NB�A�Q��^������E 3��ڜ��bi��m���=��/� �%��9������V�bN$ީ�#c<��0���ĭB/Q���F~���ݤ��	[���"� P�^he�F���H��6?4yM�e�	�Ϟ�ŚV��s�\*]��=�J��(L�U*꺟�G�D�:i��d����ױ�?�#-��Au@.(;%��l<���+��/��Μ:8�O���A��_۹��X��"�GaĥuWXvd��C�&o�U�����ņ��
�2 t�u3��C��RhN�F*��绯sJs�O����4:�V�5���Ϡ�V�!DXW�����E�+�K�N!*P0��m�c\�L�4Lm�����t�jǶ�S�)/�պ�)<� �l�|W1�]�>Gb��/�d)V46�Et������g��/%%��j��YrUh����_�pU`�.����6H�6�ަ��;�-�
�){`��~�V����rd���IS^Po�'���F�9�Hwg�Jj�{b�2A��Q�k��@O����t���������8.��~}��� d����i�e�K�L�??K�"U�4����Mo�h
V���"5�?��
���=���`��jJ���N��~΂(��1	��|��~ E���1��l�${�.^?�O�3o��ODU�X�PY��}:��)���}qJŽ�GF�+)����8�2�%E��'�~��<+�����HX�b^�Uن#_�cr붠Y+5��ޘ%��K�h1T�5��{�<RW_/l���~E�����q~�k�-p��C��{7s���8�M��SPm��*lg�A�j�,�
W)V�����:;�Ì��U#̢�,$�y� '�䗘�;���(�NI��  %A%
�;xX����ed��qG��&!�Ο�)Az�z�[{���ɢ4�!�h���xw'!;���"�,�Ib{�2�3 �'��9T�~?���*x��F´"��h-���m|?�^����.Qи���Zb������l�}��P��l��;Ȝ�bx+J�-i�1�m���B����0 @�iW�A��L�b��!@�ȊfCgN����5&�H�}���d�OE8a��cEkZ��O�Sz�~�ќe�T#���)���$@[�<�BZLT�dTC����_;jA{�E�+0�|�y;�e\0�?�fo���w�P���m�dN9����u���f�����n݈>���Lڹ�8���">�i�9jh��_dT�8���3�-����eck6�|��;O��#*�L溘E&��i�����)�z��g�Q�tef��Ό &�@5��ˆ�|�8��qg`��n��8��yJ�@�N.�inr�5��:�		�f̪&7|��Mn�%���������聀���q#�ks��uZ~��Wׅ�ñq����?v�R���^��VV�_�pC�����m+3���l՟�!��f�	D�`d�1YV?��箟x����}�a��k�#�n#�Ø##�@�p�À�3������zf*դ�4(���boN�����XAT
���`"�[���U����>�#�J�5^eZ�L�O���JS5*t�4(�F=�3g�<�����t��_b���(�(~ķ����)r�$߲.���SR���X-�\�n?��mƌ	��cS����	7V���C�����9M�O���w���\�jS�y<��ޚ��l�'��I֧��j���u��=��L{J���V�xK�B 9��r7����s�Q%L�4��>�ء��{>�����c.�ֿÆh�$d�N9�%���?/���M���"��W�.]���Q����]K��D1��]%
@|�����LSw�&�a�������/5&��B�H)~K���߰T�;p7���J8�����D�J���m�3DIX��wZ��L�B"��l�T	�,�Gk��w��AET���ch���ȝ:�C,��l��<�v5Z�蜎������-�j�r�~�X})�P��"�ʵZ-�Q[�#ņ� �1��5���&�VW����%�#�a�~�� Sz��I3��W�}�U�a;GJ7����������U�|&��)���?�;��W��#Y���z�A�'YЉ�fQ�7�t$�H�b*Ŵ��G�u�]��9}X���ե�&�UF�T4�Ϥ�{@�"i� _�8'��%Y)�B�����Kz��'�LОoO^��xRǷ1���ʽm���6*7Q�]|�1=��Nn�¡���o�1��o��+g-���r��il�PkZ*eO�3G�T�rix6�-�<��sUP�^�	w� �Q�	�?8|�qʦ�7�jX���'8Q!unkt��"�TTq��X;�\������|������_&�V?��j�zJVx\��#�*`�A�"F�؀(�wT�U����*�8�~�a�7U�'�?�� "�r�	��.d�0ߌ\�{�����8I�o��
al���/A����c��~An����k���xO`��4�[���\��,��"�*Z��BXBw��w�f�A||�3s[髟@*�{Όt���K��=�dXy����e�EH]9�k���q��st���b˻UҨ\x2p��V������.�6Q�+�p�iSAp���y;�T�l������Rb2
�bቖ�i�*{n	�϶k�,}�<X����_�U!^���fT��I���--U����J^��mS���S!���5=f��d-hM�Jw#������;�{x�^��H��ٔXYW"ս�F�|a6�[Z��&HI;������*2��|Z��\ͤ����
�܃�`m�Q:5�cӑ!���*���V����m}�'Ӥ`jP��?�]�| ��,KG���r�6$k�/�N�B���c�HYNl�Q��5X��>	ٳA�|�͟���o��俘�=]��Z!&�)bx�u>�6�2�jGb���˙���g��W�,#��+�G���,�0p�����y�2N�Eӣ0�ta@�L�'lqh���9�Ǧ|�Du+����0+�P�C��Wp�p�� ,}���r�y�$��~�2o9g��8�m�Y���~�n�|�["f�J��6v%*�wە�P��1Y4x_��`A�ʣ��2;>֊�#�ː��!Y.(�$�#ނ���$L��}\쌾�-��R�Nh(��G���4B5�0v$9(��v1V���6$o�.5��w���B]�O0e��}�e�~���&��I��	`���r��=�Y����3}۪�h[�X}C��"A7�y�|߉�^�=��#3����-,��qP�"��%nb�݉�ߌ�1/g��h�Vu�q�S?�L�P5lBg佀&)���H�g��5cz^�����>�{~�}�|������('�³��aq4(������1��ԃ%w2wL�3�D-�"�@�q9��y�)�Dz��7E��wX�#���8�� ��!�GB~_K?5ů���T��r�=���ʕ��Y�@y�z��)}��T���Ŧ���9�"s䐌�ʼ5�G圅��Û�e:�	�ڥ#E7"�b����q�28�D> �,F��z��ǟ�ط�����s�"��P݂��4�@=�#|��DO��1Ve]Ĥ�4p�P�O��%�C�c'���9�'�W���o|]���ێo�b3�"�A�Q�d��t�c\y/�v��ϣ;��d}�X�� �ū��F�%媬1���?�*�|�`��)rӳ3��R#�c��E��������Jn���Ht�X�DLk��>2�ӽ��í�~.a@��E��֌U���9T��G]��oĦ�3y�;z�WR�����ea��J9Xy%R!�)E�d!s�b�5���ה�&��a����v�ؙ��!ƎES�����kh��K��ڎ�-S�u��� ��z�`e����� �$�S���3�ЙN6�ëʾ5U }��L~8I����ze5�}��1��l�hx(ű�� �����^H��E�B{�O���"�h���ͼ.aVNM{+��-�á'g���B}����y!b�0=��*�7m����$�K\C}] K��bR�O玁4�b$Ξ��d�k�H�%;U�������퍰pk��W�mV�@�[�QX��ƹ, A��+o�4�%��ʟ�q�<,�H�wsm
�G���"�C�	T*�2�6t7?�*��٫�R�@�6�j���>T�9�S�qmj���
ԙ��> {'XèϽ��~Ƕ����B8Sх�*�*��3���u[�n%��kYm���P��$������ߣQ��7�#�Op���	��+�q<�!�#�C�_�I{�dd�bz��&�U,@O�Dt;��>�9���Nw[x�=x����y������M��̬���r?��T���fދ�Of�"��EX�F��D����s1�)A%C׷Ez%tb0�U�`�Ý�>J�n���=G��qor)v#z[I��Ǥی;</�;e�UM��쩖�Lg���OM�^N1,yڃ�)��C��N�H��g?%�o��
�#�ٷ�:|(�ʜĪ����H�)�0���?����}�׾A�A���^��.;�\<<�MN�U�>�N�ؽ3���:=8�%��z�{<�°���+y^����l/Y�.5���(��g�����E-:�N��C�ώ�Cn��P��.S�)�^o�$�	�F�?Hi��5�%��MZ�tә�9>
B�q��W�ns.���;��k$��T#K��mǄ�O���wQO�X�w)(�8]��\�4.�w�U�ٖW��P	(ԡS��=2\̊jB�#v�:[��i6o�L����,l�7,\�,��s����v���[ٕ(E�l_�m�RdK
ul�,���7���.��߄t�����vW
�~n_4�6̚A��}6ϞƤ�[�������t4Mn{1�Z��_al���C�l;C����"�� _=�����%'�]NrQn��	gh��?7]��B>3#���Ի��ώCj|��7���l�셫�*��D�q_�\:+�Tg�*D���\"=2����9��\�ΎT��Mg�%����;���^��a��dr�O�Z'�A�}��oP��\C������s+��&����=-�h�]��!�����C��	A����E]ئd!���6�_M�v�Q1�}"
P�|�I����/8hB�"�o��A�ro#5N�����������oy�A�O��6���!}G�;�	�&�_�8�T�H��\%���z?J�F��S��]D�v`���j��q�lʤ����9[���Ĉ��2P췱����ƙ�������8˫!}�����t�"�Ӧ7�$�GE5�Xg���b����K&Â���5d��G���ը��e�d��ϼK�C�/��Ϙ�G�D���%k��;��e�"��.(����j��ʆ��ۙ��'�'��ؼ�g$�sώs�N������r����o�S�UJ��,���aR���,p��1�k	2"h��#ZƑ��y΢(oCu����g�D��ǿ^+0�U���JW��}eb����B@y�yEW\��;d�Ne��I���T�뛾9��. �'�d2���I�z꘦��M��v�'�1�<�����_/�e>N&9"��*�����3��B;��m�0�P"� ��n��,��T05�b�`��>����ΐl����l���	{�r7
�����E��H��`�r��]��e�����"�6�����$C��y{-�Y��q�
TªMi���r�U@*��l�9���;�9��oԩ�m�����H
Nć_Ycl��_�<,��B2r (��ðJAJo�F3~/��?h�Y
����Q�5�&�= zbd^���d����#2�y���E?$�2�fE�)40A�w�T��Ff���V(>VdE�b/��C|��"��ƨ���5��NЯ����z:���4T�Z��<'��jf�cz�y\U͌ gB���Ij��v���`4D&�P+��χ�(��2H������4�~A��5H�AZ.Y���ik���S4���i�hwoR#̤\��r�B1WRɋ*9������ϡ���u�X�H����){"�Qk?'�#�p��a}y��x.T��g��A,��V���S(�Pݷ������ǯ�U0���Y���S�'�ڕ��U�!q�d��J�v���
�����o�B��}?J�������P�'�V�ȩ��ڃL�dq޹ϑ�5&��U�'�ɱ�?�A�2 �5T$+8!T;Bz����RlZ+� �Ĩ�RK8�����Uޜ����`���x_�V0G�ɠJ����W�`ˠ�N>�F�ͼ�;��)utm2�5�c�o��<��bi �UN�s�%F��k�$Wϙ����7_�;Z���)�r��I��6p1q�J�N2+�6�	�P1�U�=�{*1��$'�d�Y� ��92u.�:"w�+>*�p�S�y{%�@;f�Z2��.[0(|�р�0��+4cl��t��ri�@3ɤW�}]�df�vJ"����x�
lz��B��5<�M{�fY�P�[)��<�)k��փ�g�,���"ۉV^�ӟ)���R��`E�K֔�Z+����ӏh�?� r�Z���719po{T{Q���D����@�^�I���`ய�[�V|
��Y��$�o"o}��9�o=�AO8�Z�Iԭ���#�+�!s�N���ĝ�ה�;6��й�8Vԍ��U�ZF,�0���T�����!N�i~T}r��ѓ����{2�MIR[[g����j�]�&R#��\k1*׼*T@��H_g6���D�&��.�$�g|`��ni4$\M.G+w[��S7�[��ϭS�+��PN�rI��V����~��|�3��*w���cɯ��N{��L`Ϥ�m��[H,1�]�Nwg�Q��%;�J�!,��H"�o��ڰӑڝ8�{J�q+�Zh�'�Ku�_����([����P̍�Ȼ��Ã�ڰS����ۈ��T��4�G�$���N�qNO�G,dd�}����υ� lJZ댮�����n��Mz��O	KۼZ��7r��^V_5���%�ʟc��=P���f�m�l45�H��)[-ޠ2�V��dᱷ��6=�"SM����T�H(�k�A\M�#��/Jf��T�;����hf��[�����	gm�CϠ�n���l׷U�����*����"��.,�4}��V�HU��BPC�a�.��)�S8�g����W�2Z����L�G8N�ők��vS137�')��[���u|�uí2�;��M����q���<F��f��T��+=}W}L�*ݴj���G�>�ZMSO^�������w��rt�AC��M�w�Nh= �.�Z������(��\�gʻ��$,1�!��RPa�&�y�ǡ����2�c�oj^����P�Юf�,u�!㨰��g��e����+b2C�h� ��p��)�
^IC^/*O3�|n5���]$j��>���F#,�ܧSu������~ (,P�M4�G�.C�Q��_-_��D�֒��T��c�ӏf��9K���|�2�خ��G1�;c�,p�(R p��t�ҩ;��r�����tB|��.����E\2�P���)�j*���9�j�j��Чy*�Ԁ�- v��`O�� MC����@+n4��5 g����E��8��~���f>� 	�|s�r��n� 1d��u�6��p�i�o�����h�D{�툽��(XuQ�Ŏ�>��L,R�x���'���17����vZ��C�?�H<կ���H]M�ߦ[��u�H]�����:B���]~q�5�\@���_�%X��z�S�8����P���KAj��0�k!�i~�Xe�;j��}��$Y�f�2+>��R�N��������C���ᜆ �,����پjM�tP��I������H Z�DG���|�m�2y(T�|��(�ye��x��y9I7oT�H�k�?�H�����ػ�e�)\q(�}�[aӱ��Z2���K{/ݫ��ތ���Q�uQy��Q D�#Z�� p�B7��G���R�9�Ǟ�:q^P�
��d
��4С~�q������TT�k%�L�YZ��C'-(B���Ҋ�rUp�ҶN��qJ��xU��
��~𻏊�&�,E�����4L#�J��dl,����u��(�'�s���-��C՘JR7c>���4e����L� ��1��r@���[h�%)�������CG_{�>�6�Gߺ�߾�3�v���[R��,R�C�Q����%mPƨ������GH����[�ãjK�!��A��T�6HE�ʧ.��z��a�/���\�����Bs��	���� jC��E�Q4�)bnx��G>��k}�ǿM~&w[4h��6����T�=��L����
���x�������&��M���2#3�'į�N?ԁ�Y��If�v�c'��@�R�v�	�B�Hq���3ŋ��p��@(��Y�I���-��o�#U�K��4��p$7h �jd�=d٘������Kb���4��(U�0�/|6;����Q�s�
��(�(]�	:H�F�Jua����R���;�/��G2L��� �e��*64�ٵ_ɸXESvS�|e%E3yW���cʦ�����%�����pٷÌ�+��%��b�~����t��t�ug�#�|�Q �*4]�`�	d����k;�{Bl�
?}X��oOJ�moР�0�sZ����;]!�����P�.�81���=��^j�.K%j$�r���b�d)�f&���Չ$�)�3��.�_��ý�&T���4Ԧ_e��:�3�ܖw�O���uU�L�N�XPa��s�e�#����97���bT+���5��;np<ʢ�+��p��ȑh��yN4�iQ�	����qq�`��8����mR�]Byڅ4k���no>��������L�6�҃Z'�*�`JDO������v�
�*�*!�G�S�f �ԃ��I�[�<�@~�;c��1��_R�'8�_���R�SJ I>ζP�QO�(�}�o��=Fw���k�7�E뗰u���ōA�ʪ"�Z$��З��ߐ�YCF+]�%� ����Ǭ0�~�sGi�=S��x�����b���bc��ѻl�)��+�P­	�dw6��@��T���#!q��w9�A>�e�ײ���zo��G�e� �� ��oTێĲwn�x Oo&�8�>w���A?�j�=s_Z��3Q�cc�֤E�y�֣5�`��~�G�C@w��g_t�y������o�;�Ė�=�J��=>��K�����Ic_IL��3�5��: ZH�ř���b�1�v�A�a�v]��	8W�M"aa���gh�,��ʍ	�C2���=]�6�ho�>�eJn$�{9I��괗���2꽯��Mn� |�#��%'IooR�w{���eX
&Q�V�xb7��uscw��5O��H���id�Y�`�N֬���%.˩��C`�=Z��tB���=�Z�p0�磖�C�}�Ά�6b�"���۵��(��Q=6M>�����S�\�vޯ49U@<��
k����K�:���M�{ ����I�g�
H/�Q1��2�Ѐ�״��؆�:����p�� �ԥm{#�G�yn�Dt��:�4�4��M&D�z�#��H]z����נ���K�<��-c����+؀Y�0w��g�70�ۯ?�s	���&�FR�ږ>o�Cs���qd\f>�b����k�ɷ���b{��X������Km˗�on�S����7郻���<�ȁ�Xݦ���=��E�_�/cv�)��y�6�����D��ߴ��@� dRT�_�
�j�_�q[&o����_B��÷��h�/�G"��Y>�?k[�z��˟;�&�^����}>A��A_{�=9�	?	�Nh��&�{�u^*��r�Da���Z�zտ8���9���}�h5��5TZ����&x�	��0mH��iS��ű'Z�]���+b����P����ܮS_�)��Q�g�tR�����3�<X�'`y�Џ��+�@f?�,nU�|/��+�g��vi��R�xa�>�^o�3�f��~����hE�*d��!�H��oʃk�џ�r\KT����c�}�߆wb�i޻�,��9�l+��rE�:�TzP���:�q�߽� 229���n���.��.1���C
�	1�����&8�1����U�U�#;�>�fJ�!�ؾ���ia&f�C�YZQ��8��G�E���Hy�/F�����ќ���/N��yj�LH̫�<�l�C��	��!�2I�L��,�,9Y\��m¦�i�p�ߊ�${�v}��/q�=�j������<���ڝ����%���%��� ����΃1������A[��v�c�\u�~�X�]�����mg�L�4'��*����M\���%TkR����$gMiU���#n����KGe����fЪ���a`�X0�]zfbRu��9t9(�+%�ܪ)	&d=NN��R�-ֳ+W�w4L	��9���H ��
��5gM���'�"A}R�D���(�<k�����z�l���Fq�uu!<������Ȓ�j���a+��d|�������7<��w����@�����𰯇��_#�?��گ
	mD7=m��?^[W�ٛ-���r�RxueǍbܒ�d����rǁ ��z�/ճާs�n��Ե%���#�b�b��+�Z4�g&�����e�8�᪠��P�w���|�$���Z��m`*[{4i)�zyN�g��#�;J�y���ǇٕkN
j�MqcIv-�)�0�rU8#�ɺ�hG�ik�̕2��E{��CD{ B�>��ҁ��V�#ZPxC�E���W^�!����VD�z��ۑk�t���{�˖)�� |o��T��rH�(��cY�MO��Wc����u�d�y�q������x���s�q]�G��0h���7Κ5E�����QB�Q�r{c��n��m�JjNӄr#*�=�M�N9_ٯ�F5��
�m3Ul��+� 5��|н4w�i���A �;vEmd*GǞ��� �*��A�|g��̮Rqc�&*x'O�7̻{l@Rʂ�*7(��#(��O��s�c���h����.�D�CB^C�@��si���߻N,��3߃�������f���Khm�O3���bq+������&�q�|����~��49�u�gPO����C7����1���S˕Da���Rڼ�E�HT/Cɖ���
p��5�60cu����B�������Ǘ&P`=S,%zb�p�0�q���gJ��S�����-Z����eb�҆��\���x��g��F9�aG5K��y����0�9w��~������1�į%ٵRj��}���<�ZN�A�Ѹ��'ĉ���q_+�P�7R�(B�����P�y	;�2܈(�"��w��Z-ֶ��q��]{�nz��Rfu���%�����������q�� l�fFq�`�\�����ys%�����>��Bf���r��vV�{s�ɢ��]�fme�p�{�=$0�Ec�����(hI�쿙�%;����"A2�]���������
(ς�ߥ�<�y�;a~���Ǝ���	�A��;`_2�5}�_	�t�,��SQzh��]s��F���H�
�^�wH�����GK&	��:	��&������}3M@�bU�8�s��xB�ͦ���Sd��}�U�~s�y�L��!�3qk!�(�G^���{���c(��/
'P�D�_��0&ƕ�*1&�.�}�����}P���>�XZ����$��14_�p�.Eg?0�.pX��}����4>�0��o��UD%�Vu'��,��3���Nz�V��[3�z�R_�8	[��PԔ)��F6���^R
�n�$�=��ݯq��.N�6��@	U����^��T\K�S���v�h�QleK,�{]�N�(Qj���h���������X�� �&AK:�UWC����#���ə���A��}-tH)��VVvH�	 �|+ڙ릖ڔ�g%q���H�?w�BW���X�̐)�����&��Ⴜ�d��Ԋb��b��\���H��M�d�P���l�e.Q<>���t����2�����<�Ge󾲪��8~�HG�$\�Q��W��v���Y��z�XL�Z�AҸ~p���%9�̯��8"ڞ�|<�ģL���cY~|�`�s'r~�ѱ ���kg2�z� Z�l�wI)ˢ���h��]O����Q~Np�h��qX0v3��.o~��][����tl�ͼƹ�m`6Vt�����#�L� ޼��f�T���b���"I�"?�@�w�Z�D`G �~�w	�CX�.�������g���9d�ۇ���z���U��ӐR���Yf��?�@����m��$�C�i�)��h���_:ZV�bu�~i:��Gd� �{9��C̣ 8�GeR�%ρyw��k6�9���Y��m��ϯ�tٮ�Af�mX�R2>g���R
ӌ�\�Л�3�G�����e����䤙<��6����}�f��<ş�1�;���pA���1ɬ?�����䁝��M�Yߴt�-�8A�k��Ӝ��U�莥8�<�8i��]壵�Y�����&���W'��};6�'xXTj�B�����h[���޳�J	�u��Av��:�tڻ5om�r	z=!�L��a� �N����?���g����n��}#d2��-�2�b%�[^��q�>$~�MTmBț�B>��1R��t��\�g�8z?������`D�e.(��Y%n=3���r����dkP:�Υ�)�=��Du���7�J�m�#�g�����H���k}[h��Z���G����N���=�Jk��/�Jqڤu���ٚ�.8��*���DK �h�ԉ��)��ͦ:'b*z�U��KKLS�B5/��=*c���zr "#+�sn�xh��>ٗ���A��y�����#���⠡��f��Bܞ�(�s}�,�x� ��)f�t�@�vt}|��m�X[A�T�kI���H�XC����|�{�ŌE��{�s1�Ň*�.����q�( Ԏ"p�|;Q����ҕ�� ë�UT�\�/ ۬����sL/C�sӑ?jg��0���� ��D��QJK� [M,.ZӾa��K�j��ȑ��gӴ�&tM`�'� ��EL�6
4͑�ƞ�,|��%�c;"k<����#C�W
_-}H@B����\%�u>�`ϝ��*\OWl.�1���!��r�p��Y����5yL�
�W�������������v���Bq�J�&�*�r��{��v�o,*B��9�D+�ϙ��RNv�	 a�����Bƭ�� $/��"�kO឵�>�3��Gۆ`(� @|�����Y
����%}�?v��k@f�~�Cт�K�t���$O�#����������x��R3�`�E�l���.����m
x�<z��ؓ��)83�yP�m�
G����q .�m�1aS#f��kaK����Q���~Κ�����&W�%��K�R�9���7�W�}ډu�g3)O�&�!R]�9ͮ�d"��3	�*"i�H�����Yc.o��^��l�7�j�$��"ꈒ����EGW�$�5�����>�v#�E)����1f��Fݭ�mF�rv
S�R�&_�r�N���!Y� ��0�$�B�E!=�VF�jI@S::m�'铽ԉy�� �<B���FבW�5�K
�-Q���[��wi�f�#\��c��0v7��� <�)�Q����`�;�4��e�s=Qh�aՑ�TӰ}+r&ç�eIf�i���w�랬Ü��^�/ཪ��5��]�=���i�X���Zn<=�&�&H���J��ݻ5�g��+��Q0�RK0'�l�g)U����_MRp��P�B��6!^�	��k�'@��9��A��a�I���=w�a�.׸f�qϏDU�܌>q����ˇCFj7�����t��_ŉ��cF#���$h.��>+w�7ރ`K�=�E�H�?	=���?[�_��w�4Y`�ͣ��0�n��cÁ���VE}w����³F����rJ�o���)Y^��������z����a��@�(N��2"7�\h9�zQ��������Mő^�-�z���b���Ԝ�cR��[�?Oh:$�ci?��+�n1���!�;&�*s(���#˜M%w���g܈3��v��j$����=�S�����L��GKVi�u='����F8��Ʊj��&,��1�&��9�!����A���{۫��P��g��J�k�T}�G���Fp�`��;R�^~b�}���	��B�W߉)����-O����Mȳ,Ba$�>�����4��Y�Ȃ�u:|��g�P�\y��m59,��d�&y9́k?Z����D��w06�֣2Ϊb:$p!&�⏍�M_E9Ч��Xڰ������}�`�V��~��!��;#����~����F�]v����@P�q�T�t>�
�!@�V�mH�\�LM���9��*ĴϺS�+_滚$%��N��{ĵ	��8-Q��fw��GZ*�������>c���P�xR%�EJ�m�5���8~�}{��Q�({��s&q3J�ʬ�r�ϔx�q��B����TIpғ�������bs���D���r*���U0d1�0s_F�l�?T�)~��ï���a�ϝ��,$�$�P��	�0G=�οe^�ݭ�D�&�~:X���Dk���"�"�CG���{K��ۊi�͌�^Y	[�c�����d�s�I����])��K�K������T&��V%����������6R���Ǖ%���v��
���ݻ�ۜ��
YΖQ��,!9V)��wc5 �L�a�g��p��!t�?������!�]=ø�v{�Pg�q�F��Q)��o�T���c��� 8��ۮ.Md<+������8�b6f��I�!��z>����/�k�yddf�"����N� ��"�f�9�S��H�~|,�� }�x���	���Qt�B*��t����L���o�t��ˢ��Ʀ,m-���`�����=VS �4�ϡ>q�cyO���h4��)U�v�&]2�����WM���B� 3+�+%�����L�ч~o �ɽ�|l�޵�#`F�&�ff�W�*`��l�1X�A{�6�h�3���q�D�(;�˺g���e��O�FA�F��|1~�̳G@��<֨���ޔ�ΐˍr�֑oPm���U��߆�L�
�����~�,v����:�.k�~c�!>]��"��Bs�%9�W-��Bw-Bzl�~\#�|��(U9���j��'�c��"e�d�m  �t[�-��F/�$�Ǳ�Y��?G,���}'|~0G�2θ��^AK�c���B?)3�͉�2�"퐼,�4W�3���i��1�~~��² fq|���u����`v�/i����" ����O�7��}Y1�*��Mi��x�TK���9���?j���dϧu��8���tvZ)�b�J`����"u! ۵��\7�M1{���y{O�+�h�r[=���>"uF��\ۉ�<���eGflk����?�*)�x��\^`gD� o�
4���?�0�8�k��>�Ef�w�A�Hy�J�����Q�Y�Š�zp5�:����YX�;��SA��	��Ŀ��LnO4���]&.�����&�R�	dF�[҃5?��(�#�h�h$ylr��yz�M^Յ�Ug�F[W�vM���8*P��p�>/��m=V����7S9�����$ϡ�����}as����!&5�N�i���i��g�10��"z����<4Lۗo@θ�/��ϵ��ݛ6�t�Ù��������v��6����gߋ����L�����w��OD"ş-��O��cى��_���K�N8��12 �P�����.b�ʞ�`O	��6#�h���p�m���0�=��ƿ�n�¼c��
��(�}4S�˖�+�>���kE��r�L���աw n@�;���������/��.0�6���NC��#�3V;��s!6G�=�[�M�j�{�:�(t���������C��]|T�ۥ���{J�ΫT��'�)7ْ�Z�P���p�����q|���v����c,�p1l?I_��&[�s�)��dJG4>����Rǚ)���1=qkX>/_���2;�Y(����2�6�7��'rE�XO��bw0�CU���W�,� ��N��w�|���6����������g3x����V�ݗ. �Ih
�3��h(�.�	�H޺D΅'���������GҦv�u�H䩧�y�4���m�e�HD��� J�C|Km=�t��:�I���A�"�%��V��2a���l��.N C �����t�˨�oLrD�Q��~�z7�.�>�]\���Z1-&���PP�d��{]���0���>�⻁f/-��G���~�ȯ��.�tK��u�P��D���Th&���"�r~j�X���n.�kE=�����^kՔ�!@�uXKT���w�JpYN�G�q�D>l�"|�eCH��2����K����S*�4� ʕ���)Y�����q�kC/��3�Y
Q������t����_�A��ܚ�!���K��e��Z��>J>�7v������f[�:��Q*s�o9�x��M�����q)��k�CK�sS����_~������R���ARn�g����
Cl���b����|-��`�b�2�㊱W�M{(�įvYts$8����L�¨s������>�Q�M���1ٵЅ����|���>@*�-I�}�IL�WI��-`z�N�ϖ�g��v�O�ߠ�
��@0G��s�$:�Á<��J���ϓ�r��8���V"��8��xx��	���s�.�05|��6g��E��@Rf)#��8_�C��I"�υ���nv��>L��Eg����#�-��1&���Y۽��m�89���*G����	��0��=�N�ly��3��y����'�U��c�����.��H�+Q�3�r�n�B%�Zw�P�� ��	߇:C�k�	v����M�r�Ŝ��_�xcI�e�����dM�kB�!H:��k��wA#�O���t��>#��B����7X^)i���0��,�Z���E�=&(_�f{|�e�������} 2G����<���7M�᾿�&��K�S�U���I�Q�C��<��ğpبC*���;-=XL�0�~��)��k`�&���;t^.���5>8�ww�_�Z����i=�X��-wo�#�k+Ջ�zĠU`�L�@K�d�rb���I�4�� ��VeZ�!�������V=I��T/݄�FA�U��[��LV�{Q&�tvr�����.���R�m�(	Q���
ķ꿄a�f��l/A��}]�N%���R���u�^�,�#<�N���I�h�Rz)B�J��*�M;�|��>����������j����ee������A� e��D��%@S��[�A'��J�ĸ�#W��$��hHo��6�:�S����1hv6�`=�W��ar�ܧ^[Xnè.d;�C����z�f2G�0oS>�4:3oٍ�>��Bd�Z�3қ;�͍7���6�;��]�ݨ�����lC�fNۛ6	�E|�I�	���,0w�0�������#�}*�D��A
t1�'���Y|��ST��\vX��1v��A�ĩH����T��it��<G��0���Ɵ`�{2�9�V��e<e2�g�O :|��k$����#�E�����k���o\%���	���}.��@$|�?P�k���k�{�K3ο2庳���q<+����M�	�{���T
MS��v�}�r�C�
=@t�͇{oH���2�;���Gt��m�����p�F&����g���␜���u��Xx�͜�S����j���]�.�v55�`	��c�*2-�j8���ͭ�L
�H]wC�G�*z0G'����m�� �jAA�_���`�N�D&�8��>j|�F+V!�I��ʗ�*�^�"���5ՙ����5��aZ��0�4𵚰]��S,���	��t�3�_?��vM�N*)Di�1����'J���ή�	��;�D��/8BzF�[g~�t}�P��SD��\���d���E�8�����fj���]
�8�Y^��h�[��jx��E�I$=�)�iSj~8QL|�o0�=`1�yo�r���T�]2J��k@��ǛNS�Wу���?��ڄWbd�4�]k�e�Wfb�DҪ�ZF��yԲ�ŏ�@�u=���%�WDo���+��%�]�r���]��"2��3Q����b����;���D�M\�P�'{��to�S�M57m}Y�R�J��ȴ���-��R��q�lw&,�E>�[�#ow�"����]��w��B�"�����T��pב};���p���[��Ny�&Kxd���T+�Z/�pbM�d�[��66�g�]T`xξЍ��5%���z󡣹sd9{w~�8I6&S3~Jic�Ԫ5 �'�R�O�|�`'Nf��P�1S��T���)��w���' �<�0*a�qb䏍��Cr�[#������z���\���Y!�0�e '*=D��v 9�q ����[d,��X��:���tC���{0���oଛ5Śg"ų���<o�;!u6��o��>ù��������>O�m�l<������j�A�����һ�P��JN�X��[R*�j3���;b�wz�-����tإ ړP^X�:DV�#ӳ4��D�д���mU�F`da�\0��A�w��.�g����KC�����#�<�Z
�5r[_��?J�).��8.�3�����i�����L�LX�y2��kr	 ԾI�(�*�CZ4�Ŝ�p"�&�6�e�wF�W�-"GVEt�e��DL�Y�>����jK�7,�w���������v=(œ��&��Yz^�_0�����NY�c8g ؅W�CQ
�ù��v����㙚�Or
tu]���s�ͭ��<�V��/�[��P�l��z�}+���O���;]:�]G�X���A���T�{�O!Y!� o�*`*��mQE��7�F�`g���`���@�_������U8IQ��C��XĠ�|�5�� ��h�<%J+jQ���̵�Nx*%mK�s~	5�;�����0�$�a�sm��Y���B1�\]Ӣ��z�L�"���=�|����(L�Q�3*�""#���M�]2�uxNFV@
��P�vP<�>e���!�S}/TE���ڼ+(jYК�<���a��q�]kʼ�ר� y�<�)�p�NH��Ћ�˂��U��NΰS#o�ll���j���Uӹ!�~��:J|Ap�2(`5�F'D�>K>�-������Jn�We��Ol|0Ad _���,>}r����\ ˋ_B#p#��M�1F֙���[d@�Z��S���kz�P>�*B�X[I٥�e�t�2����3}�WO���y=J'_��h����Y:$P,�#_�η��֌xn�2�M�)mt�� _��������Б��be^� Ylm� ���.e,���?�����H�����D�W�gH�����Uՠ<�F&���S�D�kH�-sTK\p��Z�gV��ҥS���]����x�c�g�3�Ke�ҥ.C w�y���^1
�-��=�vT�}*��H��^�?�_�H���pOѵy���fky��ѻ��a�XuR��{�������������p�.ś	����AFMS�!��aT(�(����`����~���c̕O0�����g �����Ǣ�c��ku�N�^��Ʊ�����߲꙽�E~љ
�n1u�G%g��e�4X6�ne^�~��>���!u��A>%_�;g���]ĆF��	e�ٙ�)�u�VŢE�s��f�_Sf?�igs�U�/,4��=����Ȧ�����,�Vk��&
n:m�yU��V�"�5���7`��C�W��y̭`R���G��cB=�e�T)ⱟ������vJ5�*w�����كpr��_]Nݥ눱�Ev3�Æ:C���#�N���1������Gɩ"�D���i �C�(vZP,�+̫�WL<����M�rk�����%��,���M�ʱ�/6��
�aʩ���umjb/e�a�!���^��&5��/��$��J�æ�dA*�%Uۂ�N��$�\-����I*Nn�@�
�X���3�{��w�8�{�L{��^A�#�7��*� �s��n�`=8T����:2$��?O%CB���ELZ�ϨI� �P
�~J)�� �3N��X��(�5��\��v�tPD3֜��a]��M�\�5˞��
�WD�E�A��B�O���(^�1��Bl�����xY����#�@�����m@�$6:��,��
�T)r���3ʉ�4_U\��̓�v���+�)���� ��"'cM��L�v���W�݈c��ʬ��E*��Y������1�_|B!gGjN��>>�0\�l�1�u�#�1�e�-���\�%��a�~<�����%�6Դ+Pr��w7f�4��jv��:x?¬��D{��cX�)c�C4��ĭ��ഡ��/�N��_���Z��0<s� G�8Z����9���P 	�����U�RM������P�a~�f�`���-��� sB3���n�xkjf�*oz��-�F�y��q�	�@ߏ�M#)0�b�z���l��� 6d�I�; ,P�����\vq��6V���,d�d��p�I7Yj�����U㖝�G�j�3L;.פ�!_�%��y/�ԛ���@/Ba=�����l�6�%��qK-�v��^���m���B�U�}���$+B2�4��r׋����U<�:��>�v���Uӫ�m��y�n76m��]�}8�P
�S/��Z|ͅ��:�I�����P�6 C���,hȟdX�;'Eh�z�H�<U�N8ou���-�z�"r�"ʀ����.W|��wt����-6R���z���O %Z��.Q*�~�CI��U�uXp|�u(`!&�ڤ�M;0���4��R���5/���� Y�[����fu��~��T�b�JS��Hg�	t���۝K��u���*�.^I.��\��2��7��������j����.<?�v&��I���q���m6����+ئ�@��}H�`�em镹x�)�A�����3+ӛx:]+��$��,!7��o�*�j��7r��c?Bvjs�5.%>�s�:�@�kǨ���\���������Q�y������Q%��wr�D�5nbE%���ڗ�6fH�d��+s�l%i��M�H��ԍ����� �AGY%\�H��J2!�3�\�����Y�!�>"N��L�����gq���-�w�q�X�#oT�(_+��f�S��܇�Zr�13g^�uȩ�%��F�]Gf(���� 8��s�>G�y��Yn�@T�D^��f��8�)2�;���%e��j�ϣc=���|�ZEr��FH�h��)�y���8���E Jm�6�M�'u�?M�\�t�z��_2����\#��f���1,��"N3�7�(5�J0=rx'ߡ���G�h7�s���H-yjՀ�W��p���x���R�3H��ݫ	������_��Y-^vqh��9��:V�Wy��@�4h?�m뼖�1�Mğ'�:3g>H�AQRD��'�Y��"��TϓЬ��h�ZF|�x$:R�	J~l80A"���$�����	@��=��$
��[��4X ��ܞ�;���u9Ŕb_퓩.�"!g�'�P�k{��wL�]���&�{�����:��!������z�7�fJ�Ų����:"��zc�m0��⛍�I~�u0'��-��}�j�t��&h�(O#�ȋ�"�
�Fٟ�ǲ��?�X ��������q�mN�ʎ 퀹^�Tq:l'(��+��н�v�_�����%�x�������bYkp�FHsǩxN���-l�;�b%6i��v��*�pa�ߺ.�LQ=�|�����{���47�Xe+�	Ǥ �pU�N�����mf�a�j7����T���0w��1+G�}����m3���
�ߌ��~�O��Q4I��s���r�ш�τʗ���b^�����`a�x��^0,������nd�e���m��?&�K�)7�t���$r�y�b����8/{�� �v|E`�s�W��[kD�� U�nU%�j��x�g�d�S	H��aO�2��ө�}m�"�/�䐐H�E��9X�������hK-8*�7��L���<��ZYf�:�e*�%�Gΐ�Y��$��fr��8K!�H�@n����k�b�V?v�@,&����l6l@�qׁ�Q����� ���!,R�	�1��q�_>��G��'���,o�.�C�c�ޒ���ix �o����)�5-�_��o�X�ɷ��t����N�ki&{��ȴA�Z��Ҹ,��iSe�5�`���װS���V�nW�'�i��|���NѮ��Z�p�T�}�b�Ɖէf���X`F��\���� w�tB�<F�dR[�c�Ǩ�Y�!9u0)��r(�.��
>���
ၢ=S]d^��g�:���R�?�&�TP�"��k,�3>���{�M�Kʜ;oS"��j*�=���x�;�-�����Gj=v5�����U�����W�2(�Ә1�u�0��O��z�>��n	C㽌L^д�wp&�����t9�7 �ds�pˉ�i]��j׼�tܖ�l�$�n�����b(+�7��h{Jd4֊����B�ax��`� �~���͓��"���o�n�F>V���b,���g�e���Xr�e�D� X����"f��eϘ D�H�j���궅-u<���a]�N��[�n���x f��\?Ѱ�;�>.al�K�2-�o�P����% ����7��K%K�[�t1%��F���M�Tch�wŭ�@j�/�U �<��މ�_�zQCrR�Kaa��i���$أZ� W���㑇����K����u���GC̉� %�:z�訆��aNpQ#���ɂI�޳�=��YA��M����Ó߱�~ol�B(�J�E60s#�-o\<EY�m�5l���޾�P���9�sfg���-��IEԮp�]`����	Ľi4�"��El��I�����Kę�)ذKô��g[;ȕƳs��Z�4�	+1���=^�2�c�UKy�Un��R�g��cQ�����/����%C�$.�*��B�}�y�PF��bH�"��sdFh��C����!uݏat��	o��!M=��.���nXL�>���!Ti�M}ܛ�-#���S��p,�8Q�V4I�\�9��D�������7�y��q�Z��b�i$�z*��|~y���J��%G�+�L��g�Az��0*�g��ʬ�ZA@�~%�
1BO���^)���o��qqoxtEO����塱@�a�
���of���E�D�7�|i���e!�	ځ�_�i��v�u����L���Jd&���|$F�mG��۪E������j	@d&�0
�xՆ�S��@��XΠ�Do�M��5���T����r0A�MR":hJT���L:U F\X��u&"a�[l����L�ɂUd�ݸi0
3!2_���7�ë�pLr��f~�8�	��S8Vʨ!�BR�J@E��cP�"�@�!v�AѲ�|��B�Y��``����m��m�.��C�סrǁt_��� Dek�@��V����CU`�����d�MPu�=7��)�9,����#Å럨���=
���~�?�j��{���� ��=^�r��ݒ=Q�v��	��B�^Y+0�A-��A~.��sq9���P�;N�V��ޞh�yj��z���c.Y|��A���E���g�z�D�f�3*�����V�JS|���gmTN�����F5]�ˍM�C�.z������O���S�[����]��6a���z�
ۈQ�9��I�$�23|Yv��5y*X�~����S����}��`�ԅ���.~���9!�3~{�QfY��zG4ᏸ�6lv��g6���c%��Bu�z����Yވ�)r?.F�|�BR��W��;T��KM�V��&Y�s�0uy�B�O��;��:�P�$L���_�>b�5���6����jL�"�x���@���m�f���)X|\s/}��2�NN���	��S=����&��`��?zc�)�g>���� ;�ɥ�nN`�'Zf��m�R�P����#��,Z,ۧ�ml:k3듺��N������\RT�7�Yv:����f)�R��w��e���1f�+�;B�
���#u4��^��-���%4�f��N����S�Z� ����`K�ܚ���όCzf�a�U��,��$4�&�񬞖��{���d�r"�(�^DhF6ĊK"�r�t�r1�h�4j��,��'�/�-��/�����)Ƈ�3D�[	�M"ؘ\{J����s!�ٻ�ZtD��Xp�����\��r֛5���'&�~
�ӧL��Ǔњ�F��^�ЊQ|�tc��H��u�5��y=��Q�.��:�0�s%{����{#H��[�-��?�.N��OT�֡��x�)i ��7䡋�Q�:��%Dj���ċR�Yh� �8JX��|K��<kQ��	fUP�� �Ts<������T�E/�찮�O�ݮ<R�_v	5��s��e�k�����μ�SB(�x��v�O�5W]�Lּ�L � r���H��H6�&������/�������6�׀����<����A-��Ɩ����aL��]���MO�t�I��~wv�d/��&E�ދ���j�5�khcO���b�g;_���!�n�^����n�W�x�n%6���1����/,���
����C�Zy��bf�"��  �Eq�
D�����
���/��f���mԣOPEq=Ÿu����)�����pаZC��x#�,�/����IA ���F������Yk�~��C`�,:�aN�xlq��K�����������v%m�/�^��d`A�N<�ؿ}f!�q�<7X1gS,)`�Z�0�ޗ>���A~��2�����뎺���h0�D�}-zCq����o�Q�0����#4����*e]�R��0��f�+|r�X�T�w's���i��6<��Wc�\u\հ���#�"Z��u���ӝw���Y����7Ōs���˯��D��T;�/�{�G���qA��^U��yι~���kK�>�G�����*Crb�3(yQ��h	��tg��u���0h-�^��:�D*�>��ar��oe�3KPBVW͕�фӷ7W9�tY9���mq��h��ޮ �^����}�$c� E�,���ob��142PJ�6S��dE��~�"��c>�/v�� ��8��jVYu�-q�� ��Zׄ�4��"16<>�!J�נO�[��/�L[]:[����Bl�$jx�o��"�T�|�����ϓ���5QSD]�'7��]��0!Hm
���Dܠ��i�س�Q{/n��LFM.�
d��h���҇�������ϙ	YY��9���pJړ8����Hc��F2�ԹJ�i�._}k�w`�c��˄�+P�&�̟�� Q́~oQ�7����G�[⋳�qF,�Z9@��n�9�y�v��S�_"�ڪb�/!��K1$�B�F���p@D��`&�+N�M�P���5�޴�Y�R��㻗�٦1qwgJ�;�� bzx�>�����_��3yw���o����%F�%���I��NZO��~hG�'ҟ�1�X��-"�o�i���S��m����ҟ6����.p���cw��R������V�ZK��[m��I�Ԁ!���DT[�:���f���<�/ߡ�ε�[��Æ���=����n�q%@��~Ы�	z��p�P8G��������^���J��ߵ����T����O,"|�8��l1�n�^x�D�`Fw�E�<fO^�0W`2B}�Vg�pƩ�6����8�7_<�L���Q7��w&��V��Hl���rV���I8���d��-�U��'�uaK�j�C�I��
GJm=܅���9�ɦ�-�d���
���EU��P_�6ڦ������8�Z0X(�8��~ Y��s/6~g[������a��C����3M@,Kw�7���]��b���O5��ht�tc�9��[lxzs�C� �Y�I����+M���Q�eBh����*f�?^���T.*E���CM�d\y|_�5��P��PQH=ǝx5��nf�W{�U�:�-�:d/�yC�(0x	[��SlZ��a�r��Fц��wD����,����x0tΖ����H���8E�~IMоC>7�ZK��j9\ﴪ�jb����/%�%��˰��)�P���|�I�2���ƃQ����ve<���i,0Bx��V��/����3s��^�{}*(�!}$a����r(�ݼx��B!��OS)ȸ�^�x�/�R$W����q4@�����͐�&~
.}�_��FU����&�^�ku����=g4����+�J�]�u�?�~*�}p�0E�5(�v��A����5$^[��4��ۧĭ�ﭑ��@޺Rm�"o��&�.KM�Anv�!��o��"/�6��nՒ$�	�v��4�T�2�qg��'��i��w��>X���q
9(4Nj�Ʈf��Ωkp�(A�t[C���o?��r����C��*|.ݤ\��^���^�X����5ׅ$v*,^^��Q�v�e��l%����-L��Yz�=;���~��~�������CJ	���S�6V�@l1]�X'��ܽ	�TJX���a��E��N��"���$�$#gi�k� ��)�T�Ս/[ڧ�(]^N���W�`�'�i�oV�ɡ����P�$x�b<�����%��h�) =�5�ܱS{1��K{6
��Լ)+�'����1^%�=%��y�R�����L'�{��Gˇ�W��m�l���B�b�B{`��"j��)i{�^\@HޮKɑV�n�\T���2���<�O�x������C�b��TOo��,f��}��U6ʟ����A�=�g��~�M�׭���Mӄit~��&̥V�R�l��]���
v?��׿'Q�K�M�r���N���'��*�><P5�go4<��/w���Tz`��\�7�z)�U�}�@��҇��wB�ѭ��<���R�!��^A�]+��â"�X)�E<�Զ�%���J��i��ݞ��I�#�'y�ke�� �
Fb�^rv�7Bh����j�%�c�K�'�ςI���"5��I����$�D�ؕ�&�������wSa���m�A�n��Hٰ�V�����,��c,r���\*c�R?;���>8X� 3�_��4��=!IuH/�!�~���hU ����YS�q��
y��Eb�8�=�0�G��6ٞ@N\i���%Vs�4Zy�r���R��ۑl��6��P�e*o,\W��>��=-r�O nk���/�Qu �M�ry�J����̭�s���ȕ� �9��k�b����� }�')�O�[�E����#�ӡ�
Sa��:/Dy��D#+�~�3Zâ����:�7B5�bb�
>tH�Z`��;���Sh�ՆDI����W��[&���5eP�����R$,���^ZQ�g���O���yD�7x���h"�`���f����;��}���6~
Q�_�-ܷ	�a���j��s*U�:Į��&C�t#Vg�;s'ܰ]���9�T���c�����Z�Gl>o{��J�9��X��En���4��J��2&��.R,���²N=�O,-�������Q�zQU8B�����|^�|Ő�Q.e�ǈ�M�*��)���`/͈1%��M����b��LV�B�Ԯ�(��sm&��֊�������=��F��T��IvY^]��^}�Y�]�Y;̾���45��h��7�.���|�?�,
��{3X-���J�B���QAY���B'i�����g��}����'��z��]3���)Qز��bE�%���iw�6��-�{Y��:1��ބv��� ���*܌��N\[�ܛ{���C�V�E����O�j�+��a�AfNyJ���`h��.��=�j"f�Ud_Ֆ ����6Wu^�O��jp|R���S>40�H*���˄��l.�(dq�L�z��j]��=��҄t�z�r�ޚ
����4�D���Λ�
h(��>|���r�+t:�F.C	���J�$斋���H<M� 	F=�f�ۮ��p�lV� ��B�D ,���g���rD覎��l'��]5�g�x��m�jע�k��(�0D��pݤ�����~6��5���+2�0���HUhc- ��ԭc����p_:�����O��Ŧ]YA-j�z�"m���o&���ܝ4t�B�6[7��˝ЩS#��8s��)(ѽ��#��q3��:��&�)Q7J5l���{T�cx�Ѥ�3�߱6&.�o�UD�Q醏���)�Ť�m�zF01��h�fI���F��ϲp�칱�cJIG�'����a����N�Ip��9�(��aH����m�3�cr�k���o��*���3�xւʻ�d��|>a�1���'O���󛇽����$}g�L�{A�K����ھ�oi}���O`����h� ���4K@k֛[� �<7a����¤�[Tt>���U��y�x�ڿLbaX�ć)SnDz���m�q��(� �t���%(����ae�V�_�
D�N4�HO�%v΃V�U�k's���m66To�V/�w?v�p�ދb�T2��{k�ԕ~Hj�˜o��~
�y'R���e)�<��8�ȳ3�������TBq=U�']f{���y��K�t�㡛Ce�4�#ڭi�(���u%��CӃlq���~��B�g�.6����W�K���L�m�n�pN�۸W��(�V ����f�O]�{�%dis��_ڞj\�s�H, n��LS�vX^4�F�"b��L�e$pr*�"����NT5��0�����Ec���ɲ��^�v���$|M�f����B#Y��O*&\jD�蕲��W�g�C�?�"qM3�O��Sv�$Y�a�Fh�!�=$3�8��B4�UhZ�P<[`}��T�wM��U���`�I�r0�dÞ9C�|�@Я�=�f�@q�7Å%5���U.�
�?�韓D��:����oT#�]]��7�6[�	��6܄�ō1Ҥ�TÁ��_��aث� z�=�/��� ���Y�-�ߑ�@ayj���R��^��(��u��^�`>��7�-�B
��V���'�ǐ������WQ��Vl�����zY��=�:JC
؛����N��Cz����N&���C?����n�lր���3�5��Uz�,��n�Z�_E�e��=�I�Z0��:N,r���3��xP�VO��q���(���0�E�@N���s���N� ����dP@7}��.x��lk�a���K \�s���'�q�ɺ�]\:���O���و6gv,	~��
�g�4��$��/�1��1d/̪�kl	��X���|ꕪM_�&kx�A�#|�R�WYSi'.�������3�.���N���h	'��z+�����_�Iy��)���;^�쇏'Kj��m�iP�����!i��w�

UF��	{A���LWkhó����� sYu�!��R\��.8��%^�g(�{���:�U�^�����]�~����k���?!/-}� Bq]|�v��[Y�t'�m/X�*u���Z��s
��V=�q'S}T�IW��y0�����fg�*U޵���@�����"	��<n]0N��[�#%�~d�"�qO������,<��3����r�i��h�,��|�o�J!�=�ë���	ڇm&����)���g���5r�k*�iu�Ք� ~�#�/��P�L�f����̝4��� ��x��ñ�ռ׎����Y|:ä(����3o�y� �;��̝����x9��\��#>t�9��eɭV@s/p���(�챞64��:T�Ҵީ�lJ��Ca�!�.�[�?�:�gtde01��:������j�v��DS��s�'g/�h"�X����zBԜ.U���D��=�����ht&�߱ @���"h�yX�ǚ�g�@���͡��c�H᪦�]ΰ����>�*�w���1P�VԡOh2&���?N��̣�(7��D�h�{.��H�
9��:[8�!��Q���B]0�bU�M7�)|�N�u>(X0X�K�O���7�|Tz��O��o#Xc��' AZ��ҁᄝY�V_�R���ۘ_��n�s9.54v䘲�W!�x�ȤW��N=1>�4"�����m�)��Us(�Q��se��\h��^f�@�<{���խˢ͢:�a�$.]�;�% ��v�a^�`��mw���o�E�Ը��]�ikmGly�t���j�D)r��lM������8;�DM����s�� ^َjz�z��1;s�{  ̚Dv*L�J�Xݔ�,����R]('ػ�;�����6Ԥ�X��h"M�ڦM��nm�4��3���-�2�`�Π���M���>�O��v�'��M8l�K9%;�4�P2��r�m������g�|��<�kk�&��/���YZHK^5��︉Uv��z��d@�L�ƿ=K�������C�	�z�\���I��nY��&�"��M��i�k�q[ӄ��L�X��5����H�v��dw��Gg����A���{&����J��1�ht�I�bvi~�]xδ�J��u��࠶��� M}Y�'��0��&N�/B��*߮�����.���:e���CAF��F���(H��o����0�=�1�h��PU3u&m��t�$1�+|I�A��Ҡ�P]�4��ׄ!8����G��;k�w4��Ⱥ����\�W�x�Rx�_�Q�;�ltA�kS_$b ����!�0^�oY�&�;
���7eT$�VW^Y	�B,@I�
t#Td���Z.4Q!8,6��,�y��c��Eᣒ���,_�Y#��s� �J�� �9��T�EX�vݙ���3벂A�����)�k'dmc�8��� #ĳH	h��&<V��;�}m�%Zƨ��I+����0l9���x_g�8..��8�_@�vAא�F�t
�7�8�N�ʕ8�׮b�0�:�}��H�Ss*.w|�[iWVl���Z����7�O\5|]x���������.e�L����<1�|7�w�aﻉ��U��-�%Ђ���h_}���r��6%t��K�5�����w��n��ȣpp��Fy��y��u=�T�gQ�g>����e���_=;�@�닳x888��}r2�JwEpumi=��i=q@��"�Ы�� �K�����yL�G�I�v��a�m�#���^�q�$�6��v�1��l�U���2��)&�dµ6��R�"�N��6�ܢ" �l���ԁV`1[��k�Z�h`���ڈ��3ɠ��r�U���$Y��>�U|^ʩ�=��@
qk���C*-GH��H�m��)M�o���R�ZI����S"+��xq�O5Rvw�9��|�q@ً.�E�~����B�y�_[31 �c�:��j4���ݪ��t�Q���C�ۘ �W�����}p�{�mG��ME����_%�^Z�6`�b)�u��C1�0��-�[�vh#(g�0�|�8��߮��zey1�5��*������7����	"ж;߼����=�_0f~� `c3|3ޏ�
v�br+�ٮ��ð6v�"�HG�e�C��ޒ �Z�a\��.k��<�(�����\��٣����L�sJqcR����r^#�o��_�T�o4�o�!�$����0ݖ�k?ȶ���P��v��Y���[�.-�0�¤��>9�� �Aj�y������MoG<�Noس�z�n���/�	���3n��`UW��
K�d��CV:.N[���r��A��+_�r˶EZ�>�[����g-�	 �f-1T��smܗe���h>Z߅L�d6� ��%�#��?�y`Qa֠M�:smt���ӹ8�L��/�U�x�}�'7=�f!>����H��J�n�Jn&���^���l�"��,��Rp
W`�~��?��j���-�ɀ����b>�~�xW���^﹎l�?:���Rh��	�&
m�����B�B5�{icu�x5�6#�S"��+~l�t�O�e�gn���F����!
`�N�g~t��Ӹ�d��0	�$�@i� _��'4����!T�/�ԥFA
�k�Q(t�������6}�̦��N�	�]�b���1������?
�|!�"��'��gt�^����F�: g�����WS�V�{,Lx;:�7���;�E��gz�"��]})Z	;R�Y�!��]WO��6���Qm�J:f\��<m�iW�n�<�=����ӭ���'�W����+�B�m����ǥ,�e��3�uc���t��"=�&�����bɺ�m���i�=���Z���w�"Arq���LM���4���k��{�O���W����#�F�A�,� ��$����!��ڥ:csoN_�1(������@$��/F�tl��'^3�m �v%8�oS�ҿfLE�P]��l�N'0ϋf�@�8#�ͯ���6<�������G���@S"���Gn)׮R	��L!z�|�]7D�i0x�5\�[����z'O���f׳�A𴠙�(&3����D�y��,�s��DNR�R�`�����{gv�?���s�!@�ƂR���DYW�q��isoX�e�˩�
D
�6d"B&����&���
'1�n
O�1�旴d�xx\<6����C�>P�Ӊ@�!5F��8N���n����/��ؔC7���z��V~�x�Uo�'��\�L�u��ͳd���8�fɬ�kp}ދ��+�W�X;��<nw���3.��	<)G�yy���U�� ��h֥�z��3��k]����Y���!�n���M�t3�������w0^��tD[������ʥ��@yh��}c���'�ེR�t�e�.�ށM��|��$i�6e��u�����v�=��?��lVMWߣ��Kd]��7��=��x�t5��V����*"M
1w&m4���!c�Q&b�Y1؄��!P�4mX���
D@G�D���+�s�Ɲ�d��b�Mg �PY���o�U'ڻⲬ� >��"F��m�3��!��tAzRBIQ��
�޽�|�	2�4��m�������(TF>y��ye}�0�H3�'ϿA��<���_m�=�>����ߔ8��,6�&���A�OF��e<)C���<�K�ε�<�GJ���P�F��4�sn�����TŌ9
�|\�{����4x�$�_XW�߫I/�{�/�s�s`ŀ�p�~��g��U�W�_�������h���1s.�{4>��-�G��d��%1�2����~�6�i�q�!jGȧJki�����}��o֢Ƅ�<uO����Pf�E�h3ꋎ��@�� X�_p/�M��j�Y&ۗV4+7���k7�<�R�R�k�J}
��GFP��k�H_Z��V�DF8ˇL���<��^q�ӑd�'���&W=�6@_��ҏ��܄gH!�gi��;ؽq���lB�Lk]Z)��>l$ ��AYB8ygl��q�מQ�=�Z)�w��p�puHo�}P0O-	��D~,-V9��QW=�}��IJ�^ox(�ʛQN���mM���/�<������A=�*]Z��b1!���}��V����Պ1i�~Ip�ď���REy���B������DL!G���H��:{z�T1�7��ٗ'�2��K�g�����X��P�3pk���f�.���1'���Iκf����{ͤAZ#�V���5��#��#t��bt��YS'��"���$7�Ӡ�Z�4��3��y�l�h	��a-\x3j ;�C���v�NT+g��͌��~
��4��ie/)��p+�Fy�᳤�x��t;�u�5��jq�9� Ҥ8�N�N	Ew �}{�g�J�}*�9���e1X>�a23;�e�"\�b���4E��,�V*3f=�e��@,i=�=�T='n��Jx�@�S2	�q�����"Cۨ=x>������⬤)%�3�x�>�l��j�'+���{��#�I�%���!@������*�a&��o���h�ua���&��! #��ZYn��	_rD�����T�������.{�J&� O�������u";y��j��3�z�(�d��2g�{�8�[��}l~,���{,ɦ`�.���[[�8�W���^Y,Z��]�]+�d���U��I��
�_�x�F��'��x,���uʣ��m�_�I�F���J�6~KIDb�j�@��U_�ғ��SI�4E���Bg���Y�@�*0�,���P��)��
��Be͜���I��\�A��A]�nϴ�#�����n�(��Q�~,�c�w!Eu9���q��k_ua��c�a���3 �䮤#��f�I�(V��%�@KS �L���**�ߘ	*�2�;C �T.�MRN�
$��[�d�uQ9	�EL�b�񑔢'S. �sH�v�*��ju����V�6�L�;%�a�z���N�6��
k̃�/-�#��y�%s���9$t�3J��ck|1�Qg�_����.���*"2lڛƞ���@�A
���edX��/��v*�2�j�,r`Yh� !د���w�!C��t�ވf�w�td�G% ��9G��9	��#��~E�訄��)�(6�׀b�������z��+���:��[Z�l33}�x�o�u_�����6@�	Mŧ��E��O�X�9Uv��nOD���K���l���ȝ��5t;�`O�أ򛨚�en�V�V�����q���,,`[{~��:B�_�Ov;pMˋ4��b�z�9�`��`Q9��"�C*�!Uz-�Z�O�>|x���}a��gn������j��wVޯj�i��G	�(f�K��^Q"u굨�1�4��z2E�`s[\��zpڡ�BUL]�R	�,;,DeW�v1QXG���n�'�q�H��&<�W������2oe�j$O���%s�ѿx��s��F�d��`�ė�S�$�*�X�Y8'�/nRcr�O��-� �E^�j��g�+��eG7��л��6��E("��w�`:�`���:�B��ؑT��I���lR$�jm]I=�2��2�1S�+�Ꭻ�a�xS�y�+��5
��Z��Њ��$R?�.7� �2<xl��ȫ�o����Ej��F���b2�`3#�"�ۺ�ޅ��y�� Rp=@��8��H��V��GOD�j2�R׮��������%3���~ц����]��|Y1@�G�M��� {����$ؗ�� �{�O�s34��;k��Rf���ʞ+��
3�V�"��'�$��s�R�԰:ѹ��>�x�#҃�N�$%F/�_w�\1]}�@\���;'�IVT�L<�m�����t��+����$��)���xב�p�}���Z��BVZ�ك�l��ƾ1"���<S�q���{�ڜ�����3H�9�ד�5���eO!���n�d��-�����Q�D�7�S@a�B��	m1@�s��{�	@���,��Z�%�SO�c�,#*K	^\.�$ �2�}����w��%nG�h/չ�0iI��Xv�Z
a�?��F/��1K-J�5�g()�%T�ƚ�@��~h+]n�4���(r���<��,:�Fޝ�����K��-);y<�/��[ (�sǟ�u���3�Kw֟�(�O�]v�XgOV-��YacM��1�Ȁ�,����l'�_�If*����)����5Poƥ���ޚ���J*�G,8,8�Xw����<��pYe�~hz`��놹o�Vh���X��=M�#M��F�Mn�"���ux�,�ڔ�EHFU��.�C��N?�:��а)P��y�~�����V�H/L�]��o�9h�������&ɥ:�C1�2����s@DA���K,eD�#xb�eH��S���qj_W i�<"�����=Ʀ�Q��Q�e��hJ
u�������b��-�s4��FW�H�Ϧ������	�N���Z)GI�����$%*0IR��qϫHe�P�7��9*�y��ݦ��fp���D�zX�p{��.T��2�ϠZz#n:��4�:��Ti�o��=�x�c+�Q��Ҏ{�Y�:D�?6	�в�+���l��
��42幨8���7c;@T��Z�]-�T�;�0�׶�gR��� ޲7�>/=�b0�G�O�{���2���DwO�}����~��=����������F�{���򞌝�m�\��U0�u:)���-��@��S�s#3�
�:�W�	�?�Ē��'{���"��3��C��}'�K����ڈXjN��6f@������,���xm#0Lo��i��ơ8�*&ޢ0s�SEOP��@"^�F�?��נ6%H])�~�Q���4�n�<�
�yd kv��~�U;�t;N�љٟ�l.B�Z��%\u6���Q8WU���Xh�9���"]u�[��	X�TA���,��Ҡ�����;�r��6v�W��V�ՉHB*ZW?>n4#|�y��?��k������=M�� &5S�sc�K��di)��r��I�KW	psq��G[�e�>c5�-�@�yOb�so{���l��x�/9��W!U��Og`z�C�$���K��٪�GDzUitm��.ژ9���@t�~J�Z�#8iQ��t�7���Z��f��'���U�� %���T4��#�"��5zU@1ȝS��)4_�b�j�ѭ1�P�1	]m�m�	�t��5�Ѓ�L�ȏ���}�GӁZ7�!D�{���9��A�PF��'��*���e��/-8�dPY=��Y�=<v[�'NB��!���^��s���~������ײ��މ-Uj��� &;���.��zN�B�8^�[z����Q���w�"���*O5���5ސ����wZ���ʒ�J�[x��k�93��wy	\�u�?����`TC�B��{�j%y�M��e ����Ƿ��ej_�Έ�I-0�oS���}���Y �����ۄ�����	�}�I���AS����#;4��z�Dq{�bF�oYSW{^� ��9X���]
�:Z(UG��;�V����}VRϷ_<�g��2�o�	����!S�+�m�싁>CJD��Q�c\[�$&T�U@*���)�تH�����D������{��lY�s�=
!���.�����"GԬb�_n�o�H�xTRWE"�����[��F����q"�&�ɯ���MxH¢��o,H����t�M[��׀�h\{���0�8ĸ���ڲ��=�����< h����i,�.�H�N$
�Z�9x�/�Y�x��V��Is���t���X��τ��ћK$�W{ޮ�����[m���2��V��ݱ�!h$"�{"*V�B��+���rHZ��
IN=�ݷ�+f��q�|�g�{�5J�{͟bqJ<*��w��v�� v��Y�5�v��H2s�t;$,�9@�l���~L�F�.:��HM��}`ן;�VR��v�^�Nǀ�̾�|�o���_�R2�?���A��y�MԎP�&4,�X��z\�2ӯ���ҿ|�7tB
�0k�Oy�E�Lj���-���l�� ��3�jv�hd��i~WM�o��b��߿G�z��pG�Q2&2���v����u�6�}�%�}3Bd/G���܊���S�	��~!��W���M`�������]lԗ�K\�F�CR�{��h,˦�!����X��vM*BۚK��&�~B#�n�r��m���N�����Թ� j� ��= �,�0�[�,2y#|��+�)�%.�S�PT)
npwE!$c��0ff8X��|����LF�6x�3�d�\ARIS4�)�Q�<ࠁ����Ba�6���v����)��e]@(D��FՕ����������=��؈���{�*�"�n�Gsj: ^�s����8�X��7ɾU~_�R�vn}�a��} �]B���M�'4Y88"��Q遱�<��~=��1 ����#ͷ��:N� j�S����4g�A6�����{cpɻ���[��%���#A�q��Y?P�ri&c���G2�k���*��[Z�P�Ț���L���IM$�����%�[=*j
\����Z��.���<D�b�<X��5�<�v��3���ط��� D%�#��w}�0����M��R|�5�<�%ѭ�	Z�$�ge�!7�|L��
��3��� po �pd�

t_�K&����{A��GS-��R�����c?�Z��ЀVp�σ�a�2*�J��qu����b̜&w���ڳ#	CV~�R>��3���0�r�YB��5n;�sS�&M/aw�:G�tɉ�,5L���0@ӿ_�NG���)VJG���l-����'�'������!�����o;J� �W���g"!
H)��:-KC)^O��M�S�K.�j�.%^)zC�!�UL�ٷhxҖ7�n�������"y���
�k�qՂ�/�ɜ�J��w��w�(�O�Ÿͨ��ܭ+c��UW�N�Yhh����oi%)��K'N����!t���i��{W���MC{MLo/"�B�j�[�x � ՛�{oQ��5SwӖ�~d��5\���'Ji)��d�6��2u���y�8,���]��i�O+�����QFd�1z�ܺ7�3�G9D~�o�*K�y�3
��ύ�bȭ��<���ŧ1 Žy��V��1��j�Z�]��:3�\rF��Y5��yS	��ŒFlz��Ô'�f�Y�D�J>
��n��MK ġm���a�̐AE�m:Ҋt�j�:�?"�q%��Q�q圲]h"�,�0�R�-5Q:�����u�zع!�
g����&�H�:rb������TF80KZ:���`�{��7:����ND&��_�#c���n��(<R�(	����s!���T�ќF�é���PD�נ���?� ޹�Y��lГ��ƒ<%?���I� �u]�ʞ��dg�aƴ2��� ���a���E/�7������"�D=C��8ܚ����Ef	����5>�~��l���l�^y5�o&�o��d��"��u��眘�1�}�[���m��T����-��X�!;����:�eH�E�hD��"���7�cm}{��;��F��R*y7E���Z�X����:��|��3G�Ԓt[ ��M��-�}��{f��h�8���E�2B����~ust
�~�ɛT�������$��}Q)�9!��́���t�������&�c�����Оu�H%�qdN72$�wx�6��OM������iY�"9~3�����ӵ�{���Ρ����X�1� �q킌�����u�0�g�Ȗ���0b+�X�m����~J�ސag���dD��@��C�:n�&��Z>�.{9R��h�����O^G
�L�A߁;�Г�0��2�Y��nꎛ[��[
I)�3�㫑923%�����A���dP34�<'�M9U�{
o�۟ށ`��_�:��+�#�E�A8�D��uZ��� ���c�������7H���9��ô[Qe�r۫RC��Ί�[
��
��j~�<4�k�����{,`�P��n �!�b�ܟwh&�T�L:�&)s��+���o�pp�<�3=ϥB���� ��?�5�y�ӼO�rʢ�̸3��ks��x�%L'�+G��$F�@�p�	'(p��կwuN;��\}�&fGq�f�{QP�N��$r�&�g8Wi��X���`U�jgh�۰�UA�5�e�Ϫ�M|(N/��VG�lS1&*Y�܈�3�v���z�Q��,�DR�G��v�[�{l�I�����a��#ɐ߰J�66U�;H�]K	�(��l���U����Bs9E�P��qh��X2����g՞��aʂ�%u|$�D�>_��/�ȩi�Q���՞��J�19��7���6��v�Rhm0FL~���H�� ��T�����Д�-p��(�& �J{h�{���||�;��"�LYs�PYjH?}NJ�y�/�Ӵ:]��p�Ő�����.����odcdo���w�4�T�>��� Nϖy;M��+���~�}k(�Z�d\g\���rrSe�6��Y.p��V2�>z3q(���k�kI�˹�i�\�X��4	sͺ�T0��z��>?@&�2�tQ���kB�(�Q���;�V��E���v�%�[��A��K�JL}\�а0��������Z��D���ĠoO"}.���(�>�g�2��痩�C'F	�E��J~���Vb�k�h��t�l/�P�LNqsU#�ޞS7E����5۫�#���׍��M x+z|9��7{C'�w��z˴�?�ᩊ�����	����������Ax���3������T%�^��d	|!9�+iU�r��G�G��(��ԓ�w�F�^{d+6�L}���TN�k��:I���<���|��p�]΄(!��a�Rj���鄞ðY���౦�>/���Xl�bţ�t�*0���v[r"�/�y�����yC�wBg��]�wh�3�2�Ņ��Å�R�\�fz������q0yW�=1�@��3>���~<����S���P{e�?ol[G��l!���Ka���fH0�Y��>�c~�/��HK��"���d�S�p O���V[�j�=_�o/JV?�`���8_�X���� V���U����������*j1�S\[�(����XV��;&�/���ёZ# ��u�q��ju��}!Θ�Z��+���#��<3蝪7 O}K���vv�w�IO�rhS�<Ga��E��عK8yΨ����0=g���@�$K�x�A��<�1�u��u��v����]x6��jU��0�R]3��N���L����&�;$F����-�Q\�~�0q�-F�rA�n�B��b�7�tN��*���:8Q�2�M�]�'�
SZkRfY4���d!�܏Rl ���Qv��o�N0�1�6���X�����B� �;�Ն���R ��P�[G���;L��r@�g�༳�����|���=�l����fD�6��U��yru�pPb�M*��H�(�k����?�����D��l�0��d�)���\�*�Cͺ�Z<��Υ71�����/Z� ���O�k=_<��e8�@d��w2vL�P9Wu�Pm�+�v�7����6M�v���Qoi*q���d���,ʊo�����&0& l�Ą��C}��Ϗu@uW))��nt��&�l��͖:����T��瑊f9��˖�N�f%����wS$!�[K�!�V��..���b���^����Cǟ��=�Z�\�R�:m��<�otr@�]bY�1GՐ厚���c%��`qcn������܈JR���	��E�p鴆�\9S9�$F5�z ����۲a���G�=k:Y�|W�-��Ee߭K��z��?��L�}Lps����}.�ᾨϛ�y}*N��@Zp��@۴\xl�)}Y7�ga�� ��A}��BLx���� �F�oS�u+�����C�_�-c6�X�m)��N������@;MFX�C���=j�~Nu�]��U�_^][W��+U'Ė��5�@�0�3c��t��A][-HR����T'�fH,3�J:�G��i�jA{�U/P�6�@]��{W.�2�x�0�����7�h#�2RqM�]5�;&����6)����1!�^�&p��*�t���8�� ���@	�#o�q����+�=�o�8��u<�Z�w�6W<�bATEk	t��n)���n�cS���M:4vp�2Z�p����Jo�f�YjR�d���VwT��ܨ�ї5X5yB-�|ӪIO`�%�`ͫ/*�Fm���d�VMs���p�P[�:��b�)����(�Y�=զ�~��Z�'�M���U�����L�Ln,f�0�PQ_�~��޼EB��G�_|哆�}�E�!Xl8ݡUO
�Yj�7-^l�f����H�Q�oܡ	Z^$X�ZBrD���ǘn�\&��s���I��M�+T����<"��i~�­��2$�M�r����?�"#&C�����O�w��(�l��%��Es�wk�@��s�f]{�6���P ���U��J�H�"NP�S��?o��>�|^��E�$\��d[!���C=M����z�ވ���pǶ�=������oO��4���{��CZ��i���W��E�*_�V��6���λ����;9�i.��[�O��P����Ҷc���a���9W&����i<eFO �V%h�+��|�5 �J�����GV�a�Tވ'z�=n�K�������$5q%'�����n��̐H���<!�ּ��J�S��b�������9 ����e+�SD�.�M/��)���x5����37��t����\��C���bT����U�0�3,�����#
b\��M�L�~���Q9��9X�A�O�9�}<�i���+���=�o�P��$(��Dt��{���X�m�u#a �9��!H;9E��ӿ"&�Z��vc��C9R�*>sI��s���f�;]"�Q�W6p�p���������d��r��ȉ��8Ҷ�Wmꅿ����E�P,��:����.�����"e]�T���+�2₝^���9=Dx`hKH��_X������4��� JU~�ob��ʖ{��C+ب!	�	Y��g�yE3��w�1:v��-:0iB-��/�a�M�X��s�Z�N���!}���U����%S�h�ǚ��E���n(l;S�W8L�0���y�7�-�DD?ϋ�'�e�~�-�Y�9��\QJ�.Q���@��@���o�N?�$>ճ���z�b�c\�s.K2�̭�Y`��3L[L��vip�b?:s��sAD���%��q�X�i+�3���E_>l3`����z*�!l�`���Aw��#X�cJ���^�D,�B<d��&�[Wn�˯-�<A霎\nnc�K� <o�_�Ȓ\p#��܊��@	1�T��,O-���L�5`[j)���O��z6�_*����C����Y�X�F �(N$`F}��l��{���cQ0rH(��:�4�p��A凁��[d�w�@�M}J]2�f�N�7�\P����,qe�}�
�i���cRt�.7�{�����I�4\� ��R�33��"jX��42�J�^A�4-JZ��q��ο���՛�"sP
��^�c���c�DZ��\��5���1�=G�tbPǑ*!�Ұm�tT%χѝI�W�Zu�C���N�=��\QO�p=D)�9�<�qsڪv.^���*���{��h5o�����%o���J9�߳-�б�r�ka��SN0:am��#���0EǡA���}LͰ��E���X:-)�"�W��֐br��i7()XQ�����.gq��(c���J��Mu���Q:����ۜ[�T�1��^�H�S��uWq�6~���=�� 0�r݃Z����Nv�$�KO�yH�]�-N�ؠ����:���t���F�zG���3���4�% ������![	|�X'߅�t�r�%��h?j`Y���f��r��ʙA����UJ�U䵂�pg����O���0JW7X�o���S���O&�U�DV,�G�<�[�x���d�ƗÃ��o���*�['an�q��̍'���V�|M胥=�i7���MO�T$Q�^c*�22�#�D=#��:��̘�-dc�?o=5OYS���!#�� *ɈW�'7pn�M"?���<;�g+~[og���\���}\Z�vfX��g�1 i9��0۾h��!�;B?!z���P�:CT�CPi~��W��ֳH�.?o3h�*J�uKsr�(���n����ۃ�[��OM�4o�F:I}�'_�|�RN�)LZ�[��T�fȽ|�@W+�Y��eu^1�Sh�4p�n�V+�T"��=�A=3�~""q�?�G]��:�$��W��P|�=�PM��h��������A۳�b
��y��Q�<��!�,�5|4?D<�UNr�̱"@�$fZ���ج?6�M���ZE�I]��}�q��3���U��hu��ةf��u�����<�L\H.��v�Vi�}:X��ȵ��G(��g���{zJ���_�j�ڈp� ���(Q��.��� �$nz�G���7�>n��2 �	9 ��Ȼ��;�&�I�{Sw�$�ӂqN���v�`�(��3�fo"��mB���ߎ����˖Asl��M�������[��M���LN���i�ծ���No�o���cC�_�6�ܭ�:�SiM>�A8�_�����}�,�I�=/뻰C+��u��⾍g�����J�:����ra�Vrb{["A�(%�-׌Qa�����{A���#B~pn���
w�*bV�t����,��~��si��~�{�-f��aA�����9�sr%H%��������߀K� ��k�Q���U*ʹIΕYH��]�Ui�E�Y��'���A��4�nRx���5�%� �S�i�n)t;y��0T�(W�jG��:/��t�?NDĪ�C���t����=�Ii�Uo���wS2����įQW�(,:����рv�P68���9�����vL��b8 �-��9VN��!��$�U��(��E�k���6JG��˪&nq�&�E��>��P��=�5��������Ǌ}�o�=d>���$QT��\1[ȴ.P~�"-ːz�v���ٖ�;��ɪO��~��aX%�R�����Xs߻'C�f��l�)� �Q<�D��|�h�Nb�]�:��A��W�۩�U�K��G�l5e������
☁�C9%���%%���
El�tdcd61��p\>��H����#둺���BH� s��S��A�/e1�g�m=ڌ�)����>�k�[���?`��P�<C=����T��	߾br��OK�T�;�/��_�8��6�܁R�s�Y0��f�xfc]���<P^R�]1�d<��2�<{��R �p�;�K���˱���*E�+v�c�X���.x�{�&��6��,��M���?_d��
�R �gי��U���ͣO��X�]�@*���W�G`/���B�xV�<��B+Sn$|�/�W�W��2R���0�x��-2�|�w_VVW�������H�������ܑ������r�Ź��~��v�ص+��XV����d�RG_�b�:0#���︂{�/)�t����tQ����f�h�`H���Q,�B)+������Jo�GOF���&�c�6ӦM(�o<-F��[3s�h����-�%W�>K�:��.����@��U�z*��Z�ȋ��=�7,FD��n(``�u�x"�l^5��W�a��iqȶ�2��k7�AHm�ڷ�E��B<�=JG9�8��p�o<�{��Ĺ���-��xZ0o�X*�[_�s��[��������?�������9�������h�IŖ|hb���ړD~c1&�[.G�0�?2��qxa�*���C��_D���N�Wl틢\��	���L�DuT�x��������b�=��xz��%��(��߼�|-i�o�Ɲitʧ�^�xւ✢����z}��Fh��c��ϡ��@6(��",�?�誆��Ei�K�t-Mw���u��"��W�����yL��%.�^h?�{�ǂ��O�Ĩ�Dg�����Y�7*��˷�	��ﺜ�
�C�ӎ�먵��~͚]`r�䉁�(�/������� ,$�޶gY��8����Yd�uOv�v�#,�$׼Âs<����}TPx�zJ}&�{�	�hx�����*;�f{xpO-��yj��y�j2���מ�����tG��ްJ�F`��"�;�+�,���Z�G]��i6\��f�,K�9�}�	���]y��4վ=�^�,c�՟C�I�������B�8vi[�=8�Ԕ�9U��!}�	�/da�-)L2�,��Qn.�j��*Ѥ���o�Ã;}����]��u��AF��p�ų�ǝ�ٷ��͸�)߁4G1>a_hQ1�P|/Щ���M�S;�ŐU3�B��:P�%��8��K�%���������*��l��m����$�0�6��u����F%!寙�����Xw&�U��cF,3�иil9N&���:w:���[��W8Ԇ�e��b��v�|Ũ�e��iK�7�z�@�R-3*��a��0�m�{z�iz'y/8Ix	�sXb��p��Wk�|̊UIshj�ϒ�A�)P��Gk�)N��)�]���+Y���w�Ux��q�=kr_�O�q4j
�ʨ�޼:P���� :���n� )Ue⯭)�9T~�%�-\��芐��)�%��[f.�	Ȁ���<��'���GPK�q��d�&�[3C^��x[Ll�(j�u��G�ce+���.0{�,q��&Bi�pc���^�Sx�P�N«��P��5f�pǞ�eQ��w+Ot���T���po�@Ep%�D9�%z�d�'�o���k��BoC�P���;��⭼�S����w��C	:�s��ݸ��ßT��!f������X1Qy4x���&�q��KQW���b�|0�����k!<�c�q�$�����_x�muـ�u����2 �l����"溡�gaH`�������Ѧ"㍟����i�J. 荫�L�K��K���7�AC37N�#,+w ��L{���UH�|�����-���Q�wf�x�C��N�.s�"������\�.l�'9o~/`,QTMmhn��؊���1�{���E���aC��鹓٭���)����[�`���;�6j"�q�)?�i�(#�������%�hZT�W>����i|&�S����h�} �.'1��кpǷ]�JI��5 �wM\��ѤD��^s5�,�tvX��\�e��}Dh*�T��>��ȾbP\y h�Dc6r�b��^�-VJ���n
�����戓��_3�
�=AHזn�]�A�F%�~�����0�^�=L�����T���F#�c�H{�K���N�+ǌTz�s��C� aˍ������&�@^Jρ���7Jc���-n�������\;%-�IBk���(R8U@%���xh�l^b�`(;�gAs�	����_���C�]NS3�:�):^'��s3%�+0g$��W���{AJ�h�{�Mn+G��ە6�:s�CF=|E����s�y�,on��P��zw�xd+�{���V�.��k<����1�OZ�|������!�
��}�g���IT#i�;���7�����n�z�����HL��7Z��d�&*K���רV��"e�p��O[y�1��ӼD�@=��S��ũ�G��FdoP�p� lq�'
,Y(s3�kǅP�B/!�%��2�7�-?=L��U��������۔y{j
�~O�Aˎ:9b��&��*X�,�t��r���ⲙ�ϵ�=�=+er���6)�������M��75D~
�ѽ�;#U��=V���l�D��,Hf/ɏ_BE-��o��\eA[�y� ����ઘ9�}�z��P�w�KA�r6����;�9w 1������P�'\��Zp�/e�;1�kJ�7���L9J�	 �.�ưEN`G�3�%�x)lV�%�̅;���(-M��ّ�W�X^'�ݫ��� �<�w�m��S<Z�cY�d�D��0$�qE�&jm���л���ߛD�9o ���Cu��C��~�;Yg&�yu���dDs�MXy�c�Xp\p\�ԼSZz�d� o������*T.�a�X���:ϭ^a��B�)=��%P�Ȑ�A*۸���}��
,�B��\9�	�������%P���z$��V�y���
#1�ǋYd�ɲJ�wF�6raF�Y78�Y��d^.1`��
�{�����q�U�&���e�+C˜��jhd�U.�.��&��������DT�m�cf��aIfiӟ��`�9eFC����dK&e�����v}�"�-4���q�֓I'-j	�ξy���F,�vqE�N@���)���H�L�nuo�29j��2�l�Nׄ�c��T�?�0��AN���E��,A���7�
�s.R>+��D� �Ysv��5c�~~�]�^H.[�Ї@��A� /��N�#�L=[Z�4E��Ͽ!'̅锤_��ꖿiEG�ymX:=.�Y�^��V��_>h֯�˕2�����TV�	^���'F̷`������L�=ae"~����hh��� �;T���W�C���2<6�
��7t��ԯLZ?#S��),�ы�iF�+�3�*iʲ��'�7L��v�
[R��;�X, ���#���FIF� p��&�%=�G%=�`��58�4��څS�pΜ8��CюT�F�������I�tSé�[��4=մ��B�S����.eF���p"R=+�*�8ƶ#��I�<7n�;����Ɔ���j�U�4�<�聃�׮�;��u�Ȕ}�ҿ|;�lIX���!ې5��^�^R�.�/d+��@?2Ǡ+��:?���Q��@eW����J��R:0PY~0Snϲ�"?�x���Ǹ@��{N��YID�vJ�Jz-B�n��
��i1;ZQ\jg�`�![���/IQ!Z4�C/�M�=-i-ܭ�<T���w�d�7ʘr��e��'o:N�T5��>)MI��1�@r�ٱ:�^��6i��q��''�����Ha�{��S�����c��i����s#��?*H�&u�u�Ex`�D]<^â$��ճ}K 2�W��)[�k�d����^��W��]X,�Sʟv�
�ۉZ��o���6!��Ԁ����Ē<*�O�n�]�R�|��.?n��n����sDgm�6w�ǩ�䚚���!~`_�pk\q$�ȇ���z�$v�z��n��_!Ԥ�����{�P������s~)*N�U�HgTޚNu'5��!��O�Tp���^.3��WI�3��2�Uz��R��f�IEv�zi'q�M$����9���.���b'캈�9rA��O
��<x�k_Sx�N��x.X��}Vm��+3��G��9�����)�w`f=�����T|P�,;��dJ�
�F`���X07�n_�z�j��*�����N�A8Q9�\��H
j�v�	������$������=Jf5�;��z���[���V���"�)�#�6z�<sj,����t�Ĭ:MZ-�����ë�2&��xm�}����=��`�`����>^�W�v]yDkY�y��y�e��7g�5�S�������G�̞8�
$d\1UUy�!�C�ǿǼ�b?f�L��ĺ����kd��?�o����F�l�u(<7ǥ��N��a�
q"G�)�ZF�o�=�g�P����Yv"g�ldd�Pcv�L;Ζ7����-˯�=�ʿn[���4W�2$����5ly�ˌ0�粜.i�Q��O��!Kx�����ؖ�����垖�l����H�t���c�3~��??����]
\�]-�R>�3R��:g:�V!+�����]��1�j����N"FH�k����&�q�xl}�tֺ"h���p2A��<ud4m>;�گ��έ[�T-,U>�?�ܙ�s%�6Y��3~���P������}�Ϧ��}o�ɷ��
/��q0f��"B�w��L�I�#[����wH	��z6������&��w��=\� 	�cx4�O-��s��_�p�ϴ����V�훐���\����"�m��4�Ʈ��ץ%��T|w�Dۧ0S'��D���M��O���@ְ/+�\�#꟏�Cwɬ)�Z܂(p��ٽ{m��=H�^ tM�@q��n6� 2ŧ]�Z�ڭ}{s�2a�'��J=�CK�bx�b₣goT�;�(Hl�
