// Computer_System_camera.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System_camera (
		input  wire         alt_vip_cti_0_clocked_video_vid_clk,           //       alt_vip_cti_0_clocked_video.vid_clk
		input  wire [23:0]  alt_vip_cti_0_clocked_video_vid_data,          //                                  .vid_data
		output wire         alt_vip_cti_0_clocked_video_overflow,          //                                  .overflow
		input  wire         alt_vip_cti_0_clocked_video_vid_datavalid,     //                                  .vid_datavalid
		input  wire         alt_vip_cti_0_clocked_video_vid_locked,        //                                  .vid_locked
		input  wire         alt_vip_cti_0_clocked_video_vid_v_sync,        //                                  .vid_v_sync
		input  wire         alt_vip_cti_0_clocked_video_vid_h_sync,        //                                  .vid_h_sync
		input  wire         alt_vip_cti_0_clocked_video_vid_f,             //                                  .vid_f
		input  wire         alt_vip_vfb_0_dout_ready,                      //                alt_vip_vfb_0_dout.ready
		output wire         alt_vip_vfb_0_dout_valid,                      //                                  .valid
		output wire [23:0]  alt_vip_vfb_0_dout_data,                       //                                  .data
		output wire         alt_vip_vfb_0_dout_startofpacket,              //                                  .startofpacket
		output wire         alt_vip_vfb_0_dout_endofpacket,                //                                  .endofpacket
		input  wire         clk_clk,                                       //                               clk.clk
		input  wire [1:0]   d5m_config_avalon_av_config_slave_address,     // d5m_config_avalon_av_config_slave.address
		input  wire [3:0]   d5m_config_avalon_av_config_slave_byteenable,  //                                  .byteenable
		input  wire         d5m_config_avalon_av_config_slave_read,        //                                  .read
		input  wire         d5m_config_avalon_av_config_slave_write,       //                                  .write
		input  wire [31:0]  d5m_config_avalon_av_config_slave_writedata,   //                                  .writedata
		output wire [31:0]  d5m_config_avalon_av_config_slave_readdata,    //                                  .readdata
		output wire         d5m_config_avalon_av_config_slave_waitrequest, //                                  .waitrequest
		inout  wire         d5m_config_external_interface_SDAT,            //     d5m_config_external_interface.SDAT
		output wire         d5m_config_external_interface_SCLK,            //                                  .SCLK
		input  wire         reset_reset_n,                                 //                             reset.reset_n
		output wire [31:0]  to_ram_rd_address,                             //                         to_ram_rd.address
		output wire         to_ram_rd_read,                                //                                  .read
		input  wire         to_ram_rd_waitrequest,                         //                                  .waitrequest
		input  wire         to_ram_rd_readdatavalid,                       //                                  .readdatavalid
		input  wire [127:0] to_ram_rd_readdata,                            //                                  .readdata
		output wire [5:0]   to_ram_rd_burstcount,                          //                                  .burstcount
		output wire [31:0]  to_ram_wr_address,                             //                         to_ram_wr.address
		output wire         to_ram_wr_write,                               //                                  .write
		output wire [127:0] to_ram_wr_writedata,                           //                                  .writedata
		input  wire         to_ram_wr_waitrequest,                         //                                  .waitrequest
		output wire [3:0]   to_ram_wr_burstcount                           //                                  .burstcount
	);

	wire         alt_vip_cti_0_dout_valid;          // alt_vip_cti_0:is_valid -> alt_vip_cpr_0:din0_valid
	wire  [23:0] alt_vip_cti_0_dout_data;           // alt_vip_cti_0:is_data -> alt_vip_cpr_0:din0_data
	wire         alt_vip_cti_0_dout_ready;          // alt_vip_cpr_0:din0_ready -> alt_vip_cti_0:is_ready
	wire         alt_vip_cti_0_dout_startofpacket;  // alt_vip_cti_0:is_sop -> alt_vip_cpr_0:din0_startofpacket
	wire         alt_vip_cti_0_dout_endofpacket;    // alt_vip_cti_0:is_eop -> alt_vip_cpr_0:din0_endofpacket
	wire         alt_vip_cpr_0_dout0_valid;         // alt_vip_cpr_0:dout0_valid -> alt_vip_vfb_0:din_valid
	wire  [23:0] alt_vip_cpr_0_dout0_data;          // alt_vip_cpr_0:dout0_data -> alt_vip_vfb_0:din_data
	wire         alt_vip_cpr_0_dout0_ready;         // alt_vip_vfb_0:din_ready -> alt_vip_cpr_0:dout0_ready
	wire         alt_vip_cpr_0_dout0_startofpacket; // alt_vip_cpr_0:dout0_startofpacket -> alt_vip_vfb_0:din_startofpacket
	wire         alt_vip_cpr_0_dout0_endofpacket;   // alt_vip_cpr_0:dout0_endofpacket -> alt_vip_vfb_0:din_endofpacket

	Computer_System_camera_alt_vip_cpr_0 alt_vip_cpr_0 (
		.clock               (clk_clk),                           // clock.clk
		.reset               (~reset_reset_n),                    // reset.reset
		.din0_ready          (alt_vip_cti_0_dout_ready),          //  din0.ready
		.din0_valid          (alt_vip_cti_0_dout_valid),          //      .valid
		.din0_data           (alt_vip_cti_0_dout_data),           //      .data
		.din0_startofpacket  (alt_vip_cti_0_dout_startofpacket),  //      .startofpacket
		.din0_endofpacket    (alt_vip_cti_0_dout_endofpacket),    //      .endofpacket
		.dout0_ready         (alt_vip_cpr_0_dout0_ready),         // dout0.ready
		.dout0_valid         (alt_vip_cpr_0_dout0_valid),         //      .valid
		.dout0_data          (alt_vip_cpr_0_dout0_data),          //      .data
		.dout0_startofpacket (alt_vip_cpr_0_dout0_startofpacket), //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_0_dout0_endofpacket)    //      .endofpacket
	);

	alt_vipcti131_Vid2IS #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.SYNC_TO                       (2),
		.USE_EMBEDDED_SYNCS            (0),
		.ADD_DATA_ENABLE_SIGNAL        (0),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.USE_STD                       (0),
		.STD_WIDTH                     (1),
		.GENERATE_ANC                  (0),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS_F0            (1920),
		.V_ACTIVE_LINES_F0             (1080),
		.V_ACTIVE_LINES_F1             (32),
		.FIFO_DEPTH                    (1920),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.GENERATE_SYNC                 (0)
	) alt_vip_cti_0 (
		.is_clk        (clk_clk),                                   //       is_clk_rst.clk
		.rst           (~reset_reset_n),                            // is_clk_rst_reset.reset
		.is_data       (alt_vip_cti_0_dout_data),                   //             dout.data
		.is_valid      (alt_vip_cti_0_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_cti_0_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_cti_0_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_cti_0_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_cti_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_cti_0_clocked_video_vid_data),      //                 .export
		.overflow      (alt_vip_cti_0_clocked_video_overflow),      //                 .export
		.vid_datavalid (alt_vip_cti_0_clocked_video_vid_datavalid), //                 .export
		.vid_locked    (alt_vip_cti_0_clocked_video_vid_locked),    //                 .export
		.vid_v_sync    (alt_vip_cti_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_cti_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_cti_0_clocked_video_vid_f)          //                 .export
	);

	Computer_System_camera_alt_vip_vfb_0 alt_vip_vfb_0 (
		.clock                        (clk_clk),                           //        clock.clk
		.reset                        (~reset_reset_n),                    //        reset.reset
		.din_ready                    (alt_vip_cpr_0_dout0_ready),         //          din.ready
		.din_valid                    (alt_vip_cpr_0_dout0_valid),         //             .valid
		.din_data                     (alt_vip_cpr_0_dout0_data),          //             .data
		.din_startofpacket            (alt_vip_cpr_0_dout0_startofpacket), //             .startofpacket
		.din_endofpacket              (alt_vip_cpr_0_dout0_endofpacket),   //             .endofpacket
		.dout_ready                   (alt_vip_vfb_0_dout_ready),          //         dout.ready
		.dout_valid                   (alt_vip_vfb_0_dout_valid),          //             .valid
		.dout_data                    (alt_vip_vfb_0_dout_data),           //             .data
		.dout_startofpacket           (alt_vip_vfb_0_dout_startofpacket),  //             .startofpacket
		.dout_endofpacket             (alt_vip_vfb_0_dout_endofpacket),    //             .endofpacket
		.read_master_av_address       (to_ram_rd_address),                 //  read_master.address
		.read_master_av_read          (to_ram_rd_read),                    //             .read
		.read_master_av_waitrequest   (to_ram_rd_waitrequest),             //             .waitrequest
		.read_master_av_readdatavalid (to_ram_rd_readdatavalid),           //             .readdatavalid
		.read_master_av_readdata      (to_ram_rd_readdata),                //             .readdata
		.read_master_av_burstcount    (to_ram_rd_burstcount),              //             .burstcount
		.write_master_av_address      (to_ram_wr_address),                 // write_master.address
		.write_master_av_write        (to_ram_wr_write),                   //             .write
		.write_master_av_writedata    (to_ram_wr_writedata),               //             .writedata
		.write_master_av_waitrequest  (to_ram_wr_waitrequest),             //             .waitrequest
		.write_master_av_burstcount   (to_ram_wr_burstcount)               //             .burstcount
	);

	Computer_System_camera_d5m_config d5m_config (
		.clk         (clk_clk),                                       //                    clk.clk
		.reset       (~reset_reset_n),                                //                  reset.reset
		.address     (d5m_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (d5m_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (d5m_config_avalon_av_config_slave_read),        //                       .read
		.write       (d5m_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (d5m_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (d5m_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (d5m_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (d5m_config_external_interface_SDAT),            //     external_interface.export
		.I2C_SCLK    (d5m_config_external_interface_SCLK)             //                       .export
	);

endmodule
